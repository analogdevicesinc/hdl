// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module ad_cmos_clk #(

  parameter   DEVICE_TYPE   = 0) (

  input                   rst,
  output                  locked,

  input                   clk_in,
  output                  clk);

  localparam  SERIES7       = 0;
  localparam  VIRTEX6       = 1;

  // wires

  wire      clk_ibuf_s;

  // defaults

  assign locked = 1'b1;

  // instantiations

  IBUFG i_rx_clk_ibuf (
    .I (clk_in),
    .O (clk_ibuf_s));

  generate
  if (DEVICE_TYPE == VIRTEX6) begin
  BUFR #(.BUFR_DIVIDE("BYPASS")) i_clk_rbuf (
    .CLR (1'b0),
    .CE (1'b1),
    .I (clk_ibuf_s),
    .O (clk));
  end else begin
  BUFG i_clk_gbuf (
    .I (clk_ibuf_s),
    .O (clk));
  end
  endgenerate

endmodule

// ***************************************************************************
// ***************************************************************************

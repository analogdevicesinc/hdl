// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module axi_ad7616_maxis2wrfifo #(

  parameter   DATA_WIDTH = 16) (

  input                   clk,
  input                   rstn,
  input                   sync_in,

  // m_axis interface

  input       [DATA_WIDTH-1:0]  m_axis_data,
  output  reg             m_axis_ready,
  input                   m_axis_valid,
  output  reg             m_axis_xfer_req,

  // write fifo interface

  output  reg             fifo_wr_en,
  output  reg [DATA_WIDTH-1:0]  fifo_wr_data,
  output  reg             fifo_wr_sync,
  input                   fifo_wr_xfer_req
);


  always @(posedge clk) begin
    if (rstn == 1'b0) begin
      m_axis_ready <= 1'b0;
      m_axis_xfer_req <= 1'b0;
      fifo_wr_data <= 'b0;
      fifo_wr_en <= 1'b0;
      fifo_wr_sync <= 1'b0;
    end else begin
      m_axis_ready <= 1'b1;
      m_axis_xfer_req <= fifo_wr_xfer_req;
      fifo_wr_data <= m_axis_data;
      fifo_wr_en <= m_axis_valid;
      if (sync_in == 1'b1) begin
        fifo_wr_sync <= 1'b1;
      end else if ((m_axis_valid == 1'b1) &&
                   (fifo_wr_sync == 1'b1)) begin
        fifo_wr_sync <= 1'b0;
      end
    end
  end

endmodule

// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module fmcomms11_spi (

  // 4 wire

  input   [ 2:0]  spi_csn,
  input           spi_clk,
  input           spi_mosi,
  output          spi_miso,

  // 3 wire

  output          spi_csn_ad9625,
  output          spi_csn_ad9162,
  output          spi_csn_ad9508,
  output          spi_csn_adl5240,
  output          spi_csn_adf4355,
  output          spi_csn_hmc1119,
  inout           spi_sdio,
  output          spi_dir);

  // internal registers

  reg     [ 5:0]  spi_count = 'd0;
  reg             spi_rd_wr_n = 'd0;
  reg             spi_enable = 'd0;

  // internal signals

  wire    [ 5:0]  spi_csn6_s;
  wire            spi_csn_s;
  wire            spi_enable_s;

  // check on rising edge and change on falling edge

  assign spi_csn_ad9625 = spi_csn6_s[0];
  assign spi_csn_ad9162 = spi_csn6_s[1];
  assign spi_csn_ad9508 = spi_csn6_s[2];
  assign spi_csn_adl5240 = spi_csn6_s[3];
  assign spi_csn_adf4355 = spi_csn6_s[4];
  assign spi_csn_hmc1119 = spi_csn6_s[5];

  assign spi_csn6_s[0] = (spi_csn == 3'b001) ? 1'b0 : 1'b1;
  assign spi_csn6_s[1] = (spi_csn == 3'b010) ? 1'b0 : 1'b1;
  assign spi_csn6_s[2] = (spi_csn == 3'b011) ? 1'b0 : 1'b1;
  assign spi_csn6_s[3] = (spi_csn == 3'b100) ? 1'b0 : 1'b1;
  assign spi_csn6_s[4] = (spi_csn == 3'b101) ? 1'b0 : 1'b1;
  assign spi_csn6_s[5] = (spi_csn == 3'b110) ? 1'b0 : 1'b1;

  assign spi_csn_s = & spi_csn6_s;
  assign spi_dir = ~spi_enable_s;
  assign spi_enable_s = spi_enable & ~spi_csn_s;

  always @(posedge spi_clk or posedge spi_csn_s) begin
    if (spi_csn_s == 1'b1) begin
      spi_count <= 6'd0;
      spi_rd_wr_n <= 1'd0;
    end else begin
      spi_count <= (spi_count < 6'h3f) ? spi_count + 1'b1 : spi_count;
      if (spi_count == 6'd0) begin
        spi_rd_wr_n <= spi_mosi;
      end
    end
  end

  always @(negedge spi_clk or posedge spi_csn_s) begin
    if (spi_csn_s == 1'b1) begin
      spi_enable <= 1'b0;
    end else begin
      if (spi_count == 6'd16) begin
        spi_enable <= spi_rd_wr_n;
      end
    end
  end

  // io buffer

  assign spi_miso = spi_sdio;
  assign spi_sdio = (spi_enable_s == 1'b1) ? 1'bz : spi_mosi;

endmodule

// ***************************************************************************
// ***************************************************************************

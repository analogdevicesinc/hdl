// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// This core  is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory of
//      the repository (LICENSE_GPL2), and at: <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license as noted in the top level directory, or on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/master/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module usdrx1_spi (

  input       [ 3:0]      spi_afe_csn,
  input                   spi_clk_csn,
  input                   spi_clk,
  input                   spi_mosi,
  output                  spi_miso,

  inout                   spi_afe_sdio,
  inout                   spi_clk_sdio);

  // internal registers

  reg     [ 5:0]  spi_count = 'd0;
  reg             spi_rd_wr_n = 'd0;
  reg             spi_enable = 'd0;

  // internal signals

  wire    [ 1:0]  spi_csn_3_s;
  wire            spi_csn_s;
  wire            spi_enable_s;
  wire            spi_afe_miso_s;
  wire            spi_clk_miso_s;

  // check on rising edge and change on falling edge

  assign spi_csn_3_s[1] = & spi_afe_csn;
  assign spi_csn_3_s[0] = spi_clk_csn;
  assign spi_csn_s = & spi_csn_3_s;
  assign spi_enable_s = spi_enable & ~spi_csn_s;

  always @(posedge spi_clk or posedge spi_csn_s) begin
    if (spi_csn_s == 1'b1) begin
      spi_count <= 6'd0;
      spi_rd_wr_n <= 1'd0;
    end else begin
      spi_count <= (spi_count < 6'h3f) ? spi_count + 1'b1 : spi_count;
      if (spi_count == 6'd0) begin
        spi_rd_wr_n <= spi_mosi;
      end
    end
  end

  always @(negedge spi_clk or posedge spi_csn_s) begin
    if (spi_csn_s == 1'b1) begin
      spi_enable <= 1'b0;
    end else begin
      if (((spi_count == 6'd16)  && (spi_csn_3_s[1] == 1'b0)) ||
          ((spi_count == 6'd16) && (spi_csn_3_s[0] == 1'b0))) begin
        spi_enable <= spi_rd_wr_n;
      end
    end
  end

  assign spi_miso =  ((spi_afe_miso_s  & ~spi_csn_3_s[1]) |
                      (spi_clk_miso_s  & ~spi_csn_3_s[0]));

  // io buffers

  assign spi_afe_miso_s = spi_afe_sdio;
  assign spi_afe_sdio = (spi_enable_s == 1'b1) ? 1'bz : spi_mosi;

  assign spi_clk_miso_s = spi_clk_sdio;
  assign spi_clk_sdio = (spi_enable_s == 1'b1) ? 1'bz : spi_mosi;

endmodule

// ***************************************************************************
// ***************************************************************************

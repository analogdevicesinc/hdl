`timescale 1ns / 1ps
`default_nettype none
`include "../defs/mod_bit_cmd.vh"

module rw_register_module_tb;
	logic l_reset;
	logic l_clk = 0;
	logic l_start;
	logic [7:0] l_address = 8'hff;
	logic l_terminate = 0;

	wire w_start_ready;
	wire w_scl;
	wire w_sdi;
	wire w_sdo;
	wire w_sda;
	wire w_push_pull_en;
	wire w_error;
	wire [`MOD_BIT_CMD_WIDTH:0] w_cmd;
	wire w_cmd_tick;
	wire [7:0] w_transfer;
	wire w_transfer_valid;
	wire w_transfer_last;
	wire w_clk_quarter;
	wire w_clk_quarter;

	bit [7:0] generic_address = 8'hff;

	clk_quarter dut_clk_quarter(
		.i_reset(l_reset),
		.i_clk(l_clk),
		.o_clk(w_clk_quarter)
	);

	rw_register_module dut_rw_register_module(
		.i_reset(l_reset),
		.i_clk(l_clk),
		.i_clk_quarter(w_clk_quarter),
		.i_start(l_start),
		.o_start_ready(w_start_ready),
		.i_address(l_address),
		.i_terminate(l_terminate),

		.i_sdo(w_sdo),
		.o_cmd(w_cmd),

		.o_transfer(w_transfer),
		.o_transfer_valid(w_transfer_valid),
		.o_transfer_last(w_transfer_last),

		.o_error(w_error)
	);

	mod_bit dut_mod_bit(
		.i_reset(l_reset),
		.i_clk(l_clk),
		.i_clk_quarter(w_clk_quarter),
		.i_cmd(w_cmd),
		.o_cmd_tick(w_cmd_tick),

		.o_scl(w_scl),
		.o_sdi(w_sdi),
		.o_push_pull_en(w_push_pull_en)
	);

	phy_sda dut_phy_sda(
		.o_sdo(w_sdo),
		.i_sdi(w_sdi),
		.i_push_pull_en(w_push_pull_en),

		.io_sda(w_sda)
	);

	always #2 l_clk = ~l_clk;

	`define DUT $root.rw_register_module_tb.dut_rw_register_module
	`define TASK_CLOCK_EDGE posedge `DUT.r_clk_quarter
	task acknowledge();
		begin
			`define ACKNOWLEDGE_CONDITION \
				(`DUT.r_sm == 4) || \
				(`DUT.r_sm == 7)
			forever begin // Acknowledge or seek condition
				if (`ACKNOWLEDGE_CONDITION) begin
					force w_sdo = 1'b0;
					@(`TASK_CLOCK_EDGE);
					release w_sdo;
					break;
				end else
					@(`TASK_CLOCK_EDGE);
			end
		end
	endtask

	initial begin
		l_reset = 1'b1;
		l_start = 1'b0;

		# 10
		@(posedge l_clk);
		l_reset = 1'b0;

		@(posedge l_clk);
		@(posedge l_clk);
		@(posedge l_clk);
		@(posedge l_clk);
		@(posedge l_clk);
		l_start = 1'b1;
		@(posedge l_clk);
		l_start = 1'b0;
		@(posedge l_clk);
		acknowledge(); // Required
		acknowledge(); // Required

		#300
		l_terminate = 1'b1;
		#300

		$display("Test passed.");
		$finish;
	end

endmodule

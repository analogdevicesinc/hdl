// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// This core  is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory of
//      the repository (LICENSE_GPL2), and at: <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license as noted in the top level directory, or on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/master/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module ad_rst (

  // clock reset

  input                   preset,
  input                   clk,
  output  reg             rst);

  // internal registers

  reg             ad_rst_sync_m1 = 'd0 /* synthesis preserve */;
  reg             ad_rst_sync = 'd0 /* synthesis preserve */;

  // simple reset gen

  always @(posedge clk) begin
    ad_rst_sync_m1 <= preset;
    ad_rst_sync <= ad_rst_sync_m1;
    rst <= ad_rst_sync;
  end

endmodule

// ***************************************************************************
// ***************************************************************************

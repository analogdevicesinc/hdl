// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/100ps

module m2k_spi (

  // 4-wire

  input           ad9963_csn,
  input           adf4360_cs,
  input           spi_clk,
  input           spi_mosi,
  output          spi_miso,

  // 3-wire

  inout           spi_sdio);

  // internal registers

  reg     [ 5:0]  spi_count = 'd0;
  reg             spi_rd_wr_n = 'd0;
  reg             spi_enable = 'd0;

  // check on rising edge and change on falling edge

  always @(posedge spi_clk or posedge ad9963_csn) begin
    if (ad9963_csn == 1'b1) begin
      spi_count <= 6'd0;
      spi_rd_wr_n <= 1'd0;
    end else begin
      spi_count <= spi_count + 1'b1;
      if (spi_count == 6'd0) begin
        spi_rd_wr_n <= spi_mosi;
      end
    end
  end

  always @(negedge spi_clk or posedge ad9963_csn) begin
    if (ad9963_csn == 1'b1) begin
      spi_enable <= 1'b0;
    end else begin
      if ((spi_count == 6'd16) && (ad9963_csn == 1'b0)) begin
        spi_enable <= spi_rd_wr_n;
      end
    end
  end

  // io buffers

  assign spi_miso = spi_sdio;
  assign spi_sdio = (spi_enable == 1'b1) ? 1'bz : spi_mosi;

endmodule

// ***************************************************************************
// ***************************************************************************

// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// This core  is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory of
//      the repository (LICENSE_GPL2), and at: <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license as noted in the top level directory, or on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/master/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/1ps

module util_adxcvr_xch #(

  // parameters

  parameter   integer XCVR_ID = 0,
  parameter   integer XCVR_TYPE = 0,

  parameter   integer CPLL_FBDIV = 2,
  parameter   integer CPLL_FBDIV_4_5 = 5,

  parameter   integer TX_OUT_DIV = 1,
  parameter   integer TX_CLK25_DIV = 20,

  parameter   integer RX_OUT_DIV = 1,
  parameter   integer RX_CLK25_DIV = 20,
  parameter   [15:0]  RX_DFE_LPM_CFG = 16'h0104,
  parameter   [31:0]  RX_PMA_CFG = 32'h001e7080,
  parameter   [72:0]  RX_CDR_CFG = 72'h0b000023ff10400020) (

  // pll interface

  input           qpll2ch_clk,
  input           qpll2ch_ref_clk,
  input           qpll2ch_locked,
  input           cpll_ref_clk,
  input           up_cpll_rst,

  // receive

  input           rx_p,
  input           rx_n,

  output          rx_out_clk,
  input           rx_clk,
  output  [ 3:0]  rx_charisk,
  output  [ 3:0]  rx_disperr,
  output  [ 3:0]  rx_notintable,
  output  [31:0]  rx_data,
  input           rx_calign,

  // transmit

  output          tx_p,
  output          tx_n,

  output          tx_out_clk,
  input           tx_clk,
  input   [ 3:0]  tx_charisk,
  input   [31:0]  tx_data,

  // up interface

  input           up_rstn,
  input           up_clk,
  input   [ 7:0]  up_es_sel,
  input           up_es_enb,
  input   [11:0]  up_es_addr,
  input           up_es_wr,
  input   [15:0]  up_es_wdata,
  output  [15:0]  up_es_rdata,
  output          up_es_ready,
  output          up_rx_pll_locked,
  input           up_rx_rst,
  input           up_rx_user_ready,
  output          up_rx_rst_done,
  input           up_rx_lpm_dfe_n,
  input   [ 2:0]  up_rx_rate,
  input   [ 1:0]  up_rx_sys_clk_sel,
  input   [ 2:0]  up_rx_out_clk_sel,
  input   [ 7:0]  up_rx_sel,
  input           up_rx_enb,
  input   [11:0]  up_rx_addr,
  input           up_rx_wr,
  input   [15:0]  up_rx_wdata,
  output  [15:0]  up_rx_rdata,
  output          up_rx_ready,
  output          up_tx_pll_locked,
  input           up_tx_rst,
  input           up_tx_user_ready,
  output          up_tx_rst_done,
  input           up_tx_lpm_dfe_n,
  input   [ 2:0]  up_tx_rate,
  input   [ 1:0]  up_tx_sys_clk_sel,
  input   [ 2:0]  up_tx_out_clk_sel,
  input   [ 7:0]  up_tx_sel,
  input           up_tx_enb,
  input   [11:0]  up_tx_addr,
  input           up_tx_wr,
  input   [15:0]  up_tx_wdata,
  output  [15:0]  up_tx_rdata,
  output          up_tx_ready);

  // internal registers

  reg     [15:0]  up_es_rdata_int = 'd0;
  reg             up_es_ready_int = 'd0;
  reg     [15:0]  up_rx_rdata_int = 'd0;
  reg             up_rx_ready_int = 'd0;
  reg     [15:0]  up_tx_rdata_int = 'd0;
  reg             up_tx_ready_int = 'd0;
  reg     [ 2:0]  up_sel_int = 'd0;
  reg             up_enb_int = 'd0;
  reg     [11:0]  up_addr_int = 'd0;
  reg             up_wr_int = 'd0;
  reg     [15:0]  up_wdata_int = 'd0;
  reg             up_rx_rst_done_m1 = 'd0;
  reg             up_rx_rst_done_m2 = 'd0;
  reg             up_tx_rst_done_m1 = 'd0;
  reg             up_tx_rst_done_m2 = 'd0;
  reg     [ 2:0]  rx_rate_m1 = 'd0;
  reg     [ 2:0]  rx_rate_m2 = 'd0;
  reg     [ 2:0]  tx_rate_m1 = 'd0;
  reg     [ 2:0]  tx_rate_m2 = 'd0;

  // internal signals

  wire            up_es_enb_s;
  wire            up_rx_enb_s;
  wire            up_tx_enb_s;
  wire    [15:0]  up_rdata_s;
  wire            up_ready_s;
  wire    [ 1:0]  rx_sys_clk_sel_s;
  wire            rx_out_clk_s;
  wire            rx_rst_done_s;
  wire    [ 1:0]  tx_sys_clk_sel_s;
  wire            tx_out_clk_s;
  wire            tx_rst_done_s;
  wire    [ 1:0]  rx_pll_clk_sel_s;
  wire    [ 1:0]  tx_pll_clk_sel_s;
  wire    [11:0]  rx_charisk_open_s;
  wire    [11:0]  rx_disperr_open_s;
  wire    [ 3:0]  rx_notintable_open_s;
  wire    [95:0]  rx_data_open_s;
  wire            cpll_locked_s;

  // pll

  assign up_rx_pll_locked = (up_rx_sys_clk_sel == 2'd3) ? qpll2ch_locked : cpll_locked_s;
  assign up_tx_pll_locked = (up_tx_sys_clk_sel == 2'd3) ? qpll2ch_locked : cpll_locked_s;

  // drp access

  assign up_es_rdata = up_es_rdata_int;
  assign up_es_ready = up_es_ready_int;
  assign up_rx_rdata = up_rx_rdata_int;
  assign up_rx_ready = up_rx_ready_int;
  assign up_tx_rdata = up_tx_rdata_int;
  assign up_tx_ready = up_tx_ready_int;

  assign up_es_enb_s = ((up_es_sel == XCVR_ID) ||
    (up_es_sel == 8'hff)) ? up_es_enb : 1'b0;

  assign up_rx_enb_s = ((up_rx_sel == XCVR_ID) ||
    (up_rx_sel == 8'hff)) ? up_rx_enb : 1'b0;

  assign up_tx_enb_s = ((up_tx_sel == XCVR_ID) ||
    (up_tx_sel == 8'hff)) ? up_tx_enb : 1'b0;

  always @(negedge up_rstn or posedge up_clk) begin
    if (up_rstn == 1'b0) begin
      up_es_rdata_int <= 15'd0;
      up_es_ready_int <= 1'd0;
      up_rx_rdata_int <= 15'd0;
      up_rx_ready_int <= 1'd0;
      up_tx_rdata_int <= 15'd0;
      up_tx_ready_int <= 1'd0;
      up_sel_int <= 3'd0;
      up_enb_int <= 1'd0;
      up_addr_int <= 12'd0;
      up_wr_int <= 1'd0;
      up_wdata_int <= 15'd0;
    end else begin
      if (up_sel_int == 3'b100) begin
        up_es_rdata_int <= up_rdata_s;
        up_es_ready_int <= up_ready_s;
      end else begin
        up_es_rdata_int <= 15'd0;
        up_es_ready_int <= 1'd0;
      end
      if (up_sel_int == 3'b101) begin
        up_rx_rdata_int <= up_rdata_s;
        up_rx_ready_int <= up_ready_s;
      end else begin
        up_rx_rdata_int <= 15'd0;
        up_rx_ready_int <= 1'd0;
      end
      if (up_sel_int == 3'b110) begin
        up_tx_rdata_int <= up_rdata_s;
        up_tx_ready_int <= up_ready_s;
      end else begin
        up_tx_rdata_int <= 15'd0;
        up_tx_ready_int <= 1'd0;
      end
      if (up_sel_int[2] == 1'b1) begin
        if (up_ready_s == 1'b1) begin
          up_sel_int <= 3'b000;
        end
        up_enb_int <= 1'b0;
        up_addr_int <= 12'd0;
        up_wr_int <= 1'd0;
        up_wdata_int <= 15'd0;
      end else if (up_es_enb_s == 1'b1) begin
        up_sel_int <= 3'b100;
        up_enb_int <= 1'b1;
        up_addr_int <= up_es_addr;
        up_wr_int <= up_es_wr;
        up_wdata_int <= up_es_wdata;
      end else if (up_rx_enb_s == 1'b1) begin
        up_sel_int <= 3'b101;
        up_enb_int <= 1'b1;
        up_addr_int <= up_rx_addr;
        up_wr_int <= up_rx_wr;
        up_wdata_int <= up_rx_wdata;
      end else if (up_tx_enb_s == 1'b1) begin
        up_sel_int <= 3'b110;
        up_enb_int <= 1'b1;
        up_addr_int <= up_tx_addr;
        up_wr_int <= up_tx_wr;
        up_wdata_int <= up_tx_wdata;
      end else begin
        up_sel_int <= 3'b000;
        up_enb_int <= 1'b0;
        up_addr_int <= 12'd0;
        up_wr_int <= 1'd0;
        up_wdata_int <= 15'd0;
      end
    end
  end

  assign up_rx_rst_done = up_rx_rst_done_m2;
  assign up_tx_rst_done = up_tx_rst_done_m2;

  always @(negedge up_rstn or posedge up_clk) begin
    if (up_rstn == 1'b0) begin
      up_rx_rst_done_m1 <= 'd0;
      up_rx_rst_done_m2 <= 'd0;
      up_tx_rst_done_m1 <= 'd0;
      up_tx_rst_done_m2 <= 'd0;
    end else begin
      up_rx_rst_done_m1 <= rx_rst_done_s;
      up_rx_rst_done_m2 <= up_rx_rst_done_m1;
      up_tx_rst_done_m1 <= tx_rst_done_s;
      up_tx_rst_done_m2 <= up_tx_rst_done_m1;
    end
  end

  always @(posedge rx_clk) begin
    rx_rate_m1 <= up_rx_rate;
    rx_rate_m2 <= rx_rate_m1;
  end

  always @(posedge tx_clk) begin
    tx_rate_m1 <= up_tx_rate;
    tx_rate_m2 <= tx_rate_m1;
  end

  // instantiations

  generate
  if (XCVR_TYPE == 0) begin
  BUFG i_rx_bufg (.I (rx_out_clk_s), .O (rx_out_clk));
  BUFG i_tx_bufg (.I (tx_out_clk_s), .O (tx_out_clk));
  end
  endgenerate

  generate
  if (XCVR_TYPE == 0) begin
  assign rx_sys_clk_sel_s = up_rx_sys_clk_sel;
  assign tx_sys_clk_sel_s = up_tx_sys_clk_sel;
  assign rx_pll_clk_sel_s = 2'd0;
  assign tx_pll_clk_sel_s = 2'd0;
  end
  endgenerate

  generate
  if (XCVR_TYPE == 0) begin
  GTXE2_CHANNEL #(
    .ALIGN_COMMA_DOUBLE ("FALSE"),
    .ALIGN_COMMA_ENABLE (10'b1111111111),
    .ALIGN_COMMA_WORD (4),
    .ALIGN_MCOMMA_DET ("TRUE"),
    .ALIGN_MCOMMA_VALUE (10'b1010000011),
    .ALIGN_PCOMMA_DET ("TRUE"),
    .ALIGN_PCOMMA_VALUE (10'b0101111100),
    .CBCC_DATA_SOURCE_SEL ("DECODED"),
    .CHAN_BOND_KEEP_ALIGN ("FALSE"),
    .CHAN_BOND_MAX_SKEW (1),
    .CHAN_BOND_SEQ_1_1 (10'b0000000000),
    .CHAN_BOND_SEQ_1_2 (10'b0000000000),
    .CHAN_BOND_SEQ_1_3 (10'b0000000000),
    .CHAN_BOND_SEQ_1_4 (10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_1 (10'b0000000000),
    .CHAN_BOND_SEQ_2_2 (10'b0000000000),
    .CHAN_BOND_SEQ_2_3 (10'b0000000000),
    .CHAN_BOND_SEQ_2_4 (10'b0000000000),
    .CHAN_BOND_SEQ_2_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_USE ("FALSE"),
    .CHAN_BOND_SEQ_LEN (1),
    .CLK_CORRECT_USE ("FALSE"),
    .CLK_COR_KEEP_IDLE ("FALSE"),
    .CLK_COR_MAX_LAT (12),
    .CLK_COR_MIN_LAT (8),
    .CLK_COR_PRECEDENCE ("TRUE"),
    .CLK_COR_REPEAT_WAIT (0),
    .CLK_COR_SEQ_1_1 (10'b0100000000),
    .CLK_COR_SEQ_1_2 (10'b0000000000),
    .CLK_COR_SEQ_1_3 (10'b0000000000),
    .CLK_COR_SEQ_1_4 (10'b0000000000),
    .CLK_COR_SEQ_1_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_1 (10'b0100000000),
    .CLK_COR_SEQ_2_2 (10'b0000000000),
    .CLK_COR_SEQ_2_3 (10'b0000000000),
    .CLK_COR_SEQ_2_4 (10'b0000000000),
    .CLK_COR_SEQ_2_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_USE ("FALSE"),
    .CLK_COR_SEQ_LEN (1),
    .CPLL_CFG (24'hBC07DC),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_45 (CPLL_FBDIV_4_5),
    .CPLL_INIT_CFG (24'h00001E),
    .CPLL_LOCK_CFG (16'h01E8),
    .CPLL_REFCLK_DIV (1),
    .DEC_MCOMMA_DETECT ("TRUE"),
    .DEC_PCOMMA_DETECT ("TRUE"),
    .DEC_VALID_COMMA_ONLY ("FALSE"),
    .DMONITOR_CFG (24'h000A00),
    .ES_CONTROL (6'b000000),
    .ES_ERRDET_EN ("TRUE"),
    .ES_EYE_SCAN_EN ("TRUE"),
    .ES_HORZ_OFFSET (12'h000),
    .ES_PMA_CFG (10'b0000000000),
    .ES_PRESCALE (5'b00000),
    .ES_QUALIFIER (80'h00000000000000000000),
    .ES_QUAL_MASK (80'h00000000000000000000),
    .ES_SDATA_MASK (80'h00000000000000000000),
    .ES_VERT_OFFSET (9'b000000000),
    .FTS_DESKEW_SEQ_ENABLE (4'b1111),
    .FTS_LANE_DESKEW_CFG (4'b1111),
    .FTS_LANE_DESKEW_EN ("FALSE"),
    .GEARBOX_MODE (3'b000),
    .IS_CPLLLOCKDETCLK_INVERTED (1'b0),
    .IS_DRPCLK_INVERTED (1'b0),
    .IS_GTGREFCLK_INVERTED (1'b0),
    .IS_RXUSRCLK2_INVERTED (1'b0),
    .IS_RXUSRCLK_INVERTED (1'b0),
    .IS_TXPHDLYTSTCLK_INVERTED (1'b0),
    .IS_TXUSRCLK2_INVERTED (1'b0),
    .IS_TXUSRCLK_INVERTED (1'b0),
    .OUTREFCLK_SEL_INV (2'b11),
    .PCS_PCIE_EN ("FALSE"),
    .PCS_RSVD_ATTR (48'h000000000000),
    .PD_TRANS_TIME_FROM_P2 (12'h03c),
    .PD_TRANS_TIME_NONE_P2 (8'h3c),
    .PD_TRANS_TIME_TO_P2 (8'h64),
    .PMA_RSV (RX_PMA_CFG),
    .PMA_RSV2 (16'h2050),
    .PMA_RSV3 (2'b00),
    .PMA_RSV4 (32'h00000000),
    .RXBUFRESET_TIME (5'b00001),
    .RXBUF_ADDR_MODE ("FAST"),
    .RXBUF_EIDLE_HI_CNT (4'b1000),
    .RXBUF_EIDLE_LO_CNT (4'b0000),
    .RXBUF_EN ("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE ("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN ("FALSE"),
    .RXBUF_RESET_ON_EIDLE ("FALSE"),
    .RXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .RXBUF_THRESH_OVFLW (57),
    .RXBUF_THRESH_OVRD ("TRUE"),
    .RXBUF_THRESH_UNDFLW (3),
    .RXCDRFREQRESET_TIME (5'b00001),
    .RXCDRPHRESET_TIME (5'b00001),
    .RXCDR_CFG (RX_CDR_CFG),
    .RXCDR_FR_RESET_ON_EIDLE (1'b0),
    .RXCDR_HOLD_DURING_EIDLE (1'b0),
    .RXCDR_LOCK_CFG (6'b010101),
    .RXCDR_PH_RESET_ON_EIDLE (1'b0),
    .RXDFELPMRESET_TIME (7'b0001111),
    .RXDLY_CFG (16'h001F),
    .RXDLY_LCFG (9'h030),
    .RXDLY_TAP_CFG (16'h0000),
    .RXGEARBOX_EN ("FALSE"),
    .RXISCANRESET_TIME (5'b00001),
    .RXLPM_HF_CFG (14'b00000011110000),
    .RXLPM_LF_CFG (14'b00000011110000),
    .RXOOB_CFG (7'b0000110),
    .RXOUT_DIV (RX_OUT_DIV),
    .RXPCSRESET_TIME (5'b00001),
    .RXPHDLY_CFG (24'h084020),
    .RXPH_CFG (24'h000000),
    .RXPH_MONITOR_SEL (5'b00000),
    .RXPMARESET_TIME (5'b00011),
    .RXPRBS_ERR_LOOPBACK (1'b0),
    .RXSLIDE_AUTO_WAIT (7),
    .RXSLIDE_MODE ("OFF"),
    .RX_BIAS_CFG (12'b000000000100),
    .RX_BUFFER_CFG (6'b000000),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_CLKMUX_PD (1'b1),
    .RX_CM_SEL (2'b11),
    .RX_CM_TRIM (3'b010),
    .RX_DATA_WIDTH (40),
    .RX_DDI_SEL (6'b000000),
    .RX_DEBUG_CFG (12'b000000000000),
    .RX_DEFER_RESET_BUF_EN ("TRUE"),
    .RX_DFE_GAIN_CFG (23'h020FEA),
    .RX_DFE_H2_CFG (12'b000000000000),
    .RX_DFE_H3_CFG (12'b000001000000),
    .RX_DFE_H4_CFG (11'b00011110000),
    .RX_DFE_H5_CFG (11'b00011100000),
    .RX_DFE_KL_CFG (13'b0000011111110),
    .RX_DFE_KL_CFG2 (32'h301148AC),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_DFE_LPM_HOLD_DURING_EIDLE (1'b0),
    .RX_DFE_UT_CFG (17'b10001111000000000),
    .RX_DFE_VP_CFG (17'b00011111100000011),
    .RX_DFE_XYD_CFG (13'b0000000000000),
    .RX_DISPERR_SEQ_MATCH ("TRUE"),
    .RX_INT_DATAWIDTH (1),
    .RX_OS_CFG (13'b0000010000000),
    .RX_SIG_VALID_DLY (10),
    .RX_XCLK_SEL ("RXREC"),
    .SAS_MAX_COM (64),
    .SAS_MIN_COM (36),
    .SATA_BURST_SEQ_LEN (4'b0101),
    .SATA_BURST_VAL (3'b111),
    .SATA_CPLL_CFG ("VCO_3000MHZ"),
    .SATA_EIDLE_VAL (3'b111),
    .SATA_MAX_BURST (8),
    .SATA_MAX_INIT (21),
    .SATA_MAX_WAKE (7),
    .SATA_MIN_BURST (4),
    .SATA_MIN_INIT (12),
    .SATA_MIN_WAKE (4),
    .SHOW_REALIGN_COMMA ("TRUE"),
    .SIM_CPLLREFCLK_SEL (3'b001),
    .SIM_RECEIVER_DETECT_PASS ("TRUE"),
    .SIM_RESET_SPEEDUP ("TRUE"),
    .SIM_TX_EIDLE_DRIVE_LEVEL ("X"),
    .SIM_VERSION ("4.0"),
    .TERM_RCAL_CFG (5'b10000),
    .TERM_RCAL_OVRD (1'b0),
    .TRANS_TIME_RATE (8'h0E),
    .TST_RSV (32'h00000000),
    .TXBUF_EN ("TRUE"),
    .TXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .TXDLY_CFG (16'h001F),
    .TXDLY_LCFG (9'h030),
    .TXDLY_TAP_CFG (16'h0000),
    .TXGEARBOX_EN ("FALSE"),
    .TXOUT_DIV (TX_OUT_DIV),
    .TXPCSRESET_TIME (5'b00001),
    .TXPHDLY_CFG (24'h084020),
    .TXPH_CFG (16'h0780),
    .TXPH_MONITOR_SEL (5'b00000),
    .TXPMARESET_TIME (5'b00001),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .TX_CLKMUX_PD (1'b1),
    .TX_DATA_WIDTH (40),
    .TX_DEEMPH0 (5'b00000),
    .TX_DEEMPH1 (5'b00000),
    .TX_DRIVE_MODE ("DIRECT"),
    .TX_EIDLE_ASSERT_DELAY (3'b110),
    .TX_EIDLE_DEASSERT_DELAY (3'b100),
    .TX_INT_DATAWIDTH (1),
    .TX_LOOPBACK_DRIVE_HIZ ("FALSE"),
    .TX_MAINCURSOR_SEL (1'b0),
    .TX_MARGIN_FULL_0 (7'b1001110),
    .TX_MARGIN_FULL_1 (7'b1001001),
    .TX_MARGIN_FULL_2 (7'b1000101),
    .TX_MARGIN_FULL_3 (7'b1000010),
    .TX_MARGIN_FULL_4 (7'b1000000),
    .TX_MARGIN_LOW_0 (7'b1000110),
    .TX_MARGIN_LOW_1 (7'b1000100),
    .TX_MARGIN_LOW_2 (7'b1000010),
    .TX_MARGIN_LOW_3 (7'b1000000),
    .TX_MARGIN_LOW_4 (7'b1000000),
    .TX_PREDRIVER_MODE (1'b0),
    .TX_QPI_STATUS_EN (1'b0),
    .TX_RXDETECT_CFG (14'h1832),
    .TX_RXDETECT_REF (3'b100),
    .TX_XCLK_SEL ("TXOUT"),
    .UCODEER_CLR (1'b0))
  i_gtxe2_channel (
    .RXOUTCLKPCS (),
    .RXPHSLIPMONITOR (),
    .PHYSTATUS (),
    .RXCDRLOCK (),
    .RXCHANBONDSEQ (),
    .RXCHANISALIGNED (),
    .RXCHANREALIGN (),
    .RXCOMINITDET (),
    .RXCOMSASDET (),
    .RXCOMWAKEDET (),
    .RXDATAVALID (),
    .RXDLYSRESETDONE (),
    .RXELECIDLE (),
    .RXHEADERVALID (),
    .RXPHALIGNDONE (),
    .RXQPISENN (),
    .RXQPISENP (),
    .RXRATEDONE (),
    .RXSTARTOFSEQ (),
    .RXVALID (),
    .TXCOMFINISH (),
    .TXDLYSRESETDONE (),
    .TXGEARBOXREADY (),
    .TXPHALIGNDONE (),
    .TXPHINITDONE (),
    .TXQPISENN (),
    .TXQPISENP (),
    .TXRATEDONE (),
    .PCSRSVDOUT (),
    .RXCLKCORCNT (),
    .RXHEADER (),
    .RXCHBONDO (),
    .RXPHMONITOR (),
    .TSTOUT (),
    .GTREFCLKMONITOR (),
    .CFGRESET (1'h0),
    .CLKRSVD (4'h0),
    .CPLLFBCLKLOST (),
    .CPLLLOCK (cpll_locked_s),
    .CPLLLOCKDETCLK (up_clk),
    .CPLLLOCKEN (1'h1),
    .CPLLPD (1'h0),
    .CPLLREFCLKLOST (),
    .CPLLREFCLKSEL (3'h1),
    .CPLLRESET (up_cpll_rst),
    .DMONITOROUT (),
    .DRPADDR (up_addr_int[8:0]),
    .DRPCLK (up_clk),
    .DRPDI (up_wdata_int),
    .DRPDO (up_rdata_s),
    .DRPEN (up_enb_int),
    .DRPRDY (up_ready_s),
    .DRPWE (up_wr_int),
    .EYESCANDATAERROR (),
    .EYESCANMODE (1'h0),
    .EYESCANRESET (1'h0),
    .EYESCANTRIGGER (1'h0),
    .GTGREFCLK (1'h0),
    .GTNORTHREFCLK0 (1'h0),
    .GTNORTHREFCLK1 (1'h0),
    .GTREFCLK0 (cpll_ref_clk),
    .GTREFCLK1 (1'h0),
    .GTRESETSEL (1'h0),
    .GTRSVD (16'h0),
    .GTRXRESET (up_rx_rst),
    .GTSOUTHREFCLK0 (1'h0),
    .GTSOUTHREFCLK1 (1'h0),
    .GTTXRESET (up_tx_rst),
    .GTXRXN (rx_n),
    .GTXRXP (rx_p),
    .GTXTXN (tx_n),
    .GTXTXP (tx_p),
    .LOOPBACK (3'h0),
    .PCSRSVDIN (16'h0),
    .PCSRSVDIN2 (5'h0),
    .PMARSVDIN (5'h0),
    .PMARSVDIN2 (5'h0),
    .QPLLCLK (qpll2ch_clk),
    .QPLLREFCLK (qpll2ch_ref_clk),
    .RESETOVRD (1'h0),
    .RX8B10BEN (1'h1),
    .RXBUFRESET (1'h0),
    .RXBUFSTATUS (),
    .RXBYTEISALIGNED (),
    .RXBYTEREALIGN (),
    .RXCDRFREQRESET (1'h0),
    .RXCDRHOLD (1'h0),
    .RXCDROVRDEN (1'h0),
    .RXCDRRESET (1'h0),
    .RXCDRRESETRSV (1'h0),
    .RXCHARISCOMMA (),
    .RXCHARISK ({rx_charisk_open_s[3:0], rx_charisk}),
    .RXCHBONDEN (1'h0),
    .RXCHBONDI (5'h0),
    .RXCHBONDLEVEL (3'h0),
    .RXCHBONDMASTER (1'h1),
    .RXCHBONDSLAVE (1'h0),
    .RXCOMMADET (),
    .RXCOMMADETEN (1'h1),
    .RXDATA ({rx_data_open_s[31:0], rx_data}),
    .RXDDIEN (1'h0),
    .RXDFEAGCHOLD (1'h0),
    .RXDFEAGCOVRDEN (1'h0),
    .RXDFECM1EN (1'h0),
    .RXDFELFHOLD (1'h0),
    .RXDFELFOVRDEN (1'h0),
    .RXDFELPMRESET (1'h0),
    .RXDFETAP2HOLD (1'h0),
    .RXDFETAP2OVRDEN (1'h0),
    .RXDFETAP3HOLD (1'h0),
    .RXDFETAP3OVRDEN (1'h0),
    .RXDFETAP4HOLD (1'h0),
    .RXDFETAP4OVRDEN (1'h0),
    .RXDFETAP5HOLD (1'h0),
    .RXDFETAP5OVRDEN (1'h0),
    .RXDFEUTHOLD (1'h0),
    .RXDFEUTOVRDEN (1'h0),
    .RXDFEVPHOLD (1'h0),
    .RXDFEVPOVRDEN (1'h0),
    .RXDFEVSEN (1'h0),
    .RXDFEXYDEN (1'h1),
    .RXDFEXYDHOLD (1'h0),
    .RXDFEXYDOVRDEN (1'h0),
    .RXDISPERR ({rx_disperr_open_s[3:0], rx_disperr}),
    .RXDLYBYPASS (1'h1),
    .RXDLYEN (1'h0),
    .RXDLYOVRDEN (1'h0),
    .RXDLYSRESET (1'h0),
    .RXELECIDLEMODE (2'h3),
    .RXGEARBOXSLIP (1'h0),
    .RXLPMEN (up_rx_lpm_dfe_n),
    .RXLPMHFHOLD (1'h0),
    .RXLPMHFOVRDEN (1'h0),
    .RXLPMLFHOLD (1'h0),
    .RXLPMLFKLOVRDEN (1'h0),
    .RXMCOMMAALIGNEN (rx_calign),
    .RXMONITOROUT (),
    .RXMONITORSEL (2'h0),
    .RXNOTINTABLE ({rx_notintable_open_s, rx_notintable}),
    .RXOOBRESET (1'h0),
    .RXOSHOLD (1'h0),
    .RXOSOVRDEN (1'h0),
    .RXOUTCLK (rx_out_clk_s),
    .RXOUTCLKFABRIC (),
    .RXOUTCLKSEL (up_rx_out_clk_sel),
    .RXPCOMMAALIGNEN (rx_calign),
    .RXPCSRESET (1'h0),
    .RXPD (2'h0),
    .RXPHALIGN (1'h0),
    .RXPHALIGNEN (1'h0),
    .RXPHDLYPD (1'h0),
    .RXPHDLYRESET (1'h0),
    .RXPHOVRDEN (1'h0),
    .RXPMARESET (1'h0),
    .RXPOLARITY (1'h0),
    .RXPRBSCNTRESET (1'h0),
    .RXPRBSERR (),
    .RXPRBSSEL (3'h0),
    .RXQPIEN (1'h0),
    .RXRATE (rx_rate_m2),
    .RXRESETDONE (rx_rst_done_s),
    .RXSLIDE (1'h0),
    .RXSTATUS (),
    .RXSYSCLKSEL (rx_sys_clk_sel_s),
    .RXUSERRDY (up_rx_user_ready),
    .RXUSRCLK (rx_clk),
    .RXUSRCLK2 (rx_clk),
    .SETERRSTATUS (1'h0),
    .TSTIN (20'hfffff),
    .TX8B10BBYPASS (8'h0),
    .TX8B10BEN (1'h1),
    .TXBUFDIFFCTRL (3'h4),
    .TXBUFSTATUS (),
    .TXCHARDISPMODE (8'h0),
    .TXCHARDISPVAL (8'h0),
    .TXCHARISK ({4'd0, tx_charisk}),
    .TXCOMINIT (1'h0),
    .TXCOMSAS (1'h0),
    .TXCOMWAKE (1'h0),
    .TXDATA ({32'd0, tx_data}),
    .TXDEEMPH (1'h0),
    .TXDETECTRX (1'h0),
    .TXDIFFCTRL (4'h8),
    .TXDIFFPD (1'h0),
    .TXDLYBYPASS (1'h1),
    .TXDLYEN (1'h0),
    .TXDLYHOLD (1'h0),
    .TXDLYOVRDEN (1'h0),
    .TXDLYSRESET (1'h0),
    .TXDLYUPDOWN (1'h0),
    .TXELECIDLE (1'h0),
    .TXHEADER (3'h0),
    .TXINHIBIT (1'h0),
    .TXMAINCURSOR (7'h0),
    .TXMARGIN (3'h0),
    .TXOUTCLK (tx_out_clk_s),
    .TXOUTCLKFABRIC (),
    .TXOUTCLKPCS (),
    .TXOUTCLKSEL (up_tx_out_clk_sel),
    .TXPCSRESET (1'h0),
    .TXPD (2'h0),
    .TXPDELECIDLEMODE (1'h0),
    .TXPHALIGN (1'h0),
    .TXPHALIGNEN (1'h0),
    .TXPHDLYPD (1'h0),
    .TXPHDLYRESET (1'h0),
    .TXPHDLYTSTCLK (1'h0),
    .TXPHINIT (1'h0),
    .TXPHOVRDEN (1'h0),
    .TXPISOPD (1'h0),
    .TXPMARESET (1'h0),
    .TXPOLARITY (1'h0),
    .TXPOSTCURSOR (5'h0),
    .TXPOSTCURSORINV (1'h0),
    .TXPRBSFORCEERR (1'h0),
    .TXPRBSSEL (3'd0),
    .TXPRECURSOR (5'h0),
    .TXPRECURSORINV (1'h0),
    .TXQPIBIASEN (1'h0),
    .TXQPISTRONGPDOWN (1'h0),
    .TXQPIWEAKPUP (1'h0),
    .TXRATE (tx_rate_m2),
    .TXRESETDONE (tx_rst_done_s),
    .TXSEQUENCE (7'h0),
    .TXSTARTSEQ (1'h0),
    .TXSWING (1'h0),
    .TXSYSCLKSEL (tx_sys_clk_sel_s),
    .TXUSERRDY (up_tx_user_ready),
    .TXUSRCLK (tx_clk),
    .TXUSRCLK2 (tx_clk));
  end
  endgenerate

  generate
  if (XCVR_TYPE == 1) begin
  BUFG_GT i_rx_bufg (
    .CE (1'b1),
    .CEMASK (1'b0),
    .CLR (1'b0),
    .CLRMASK (1'b0),
    .DIV (3'd0),
    .I (rx_out_clk_s),
    .O (rx_out_clk));

  BUFG_GT i_tx_bufg (
    .CE (1'b1),
    .CEMASK (1'b0),
    .CLR (1'b0),
    .CLRMASK (1'b0),
    .DIV (3'd0),
    .I (tx_out_clk_s),
    .O (tx_out_clk));
  end
  endgenerate

  generate
  if (XCVR_TYPE == 1) begin
  assign rx_sys_clk_sel_s = (up_rx_sys_clk_sel == 2'd3) ? 2'b10 : 2'b00;
  assign tx_sys_clk_sel_s = (up_tx_sys_clk_sel == 2'd3) ? 2'b10 : 2'b00;
  assign rx_pll_clk_sel_s = up_rx_sys_clk_sel;
  assign tx_pll_clk_sel_s = up_tx_sys_clk_sel;
  end
  endgenerate

  generate
  if (XCVR_TYPE == 1) begin
  GTHE3_CHANNEL #(
    .ACJTAG_DEBUG_MODE (1'b0),
    .ACJTAG_MODE (1'b0),
    .ACJTAG_RESET (1'b0),
    .ADAPT_CFG0 (16'hf800),
    .ADAPT_CFG1 (16'h0000),
    .ALIGN_COMMA_DOUBLE ("FALSE"),
    .ALIGN_COMMA_ENABLE (10'b1111111111),
    .ALIGN_COMMA_WORD (1),
    .ALIGN_MCOMMA_DET ("TRUE"),
    .ALIGN_MCOMMA_VALUE (10'b1010000011),
    .ALIGN_PCOMMA_DET ("TRUE"),
    .ALIGN_PCOMMA_VALUE (10'b0101111100),
    .A_RXOSCALRESET (1'b0),
    .A_RXPROGDIVRESET (1'b0),
    .A_TXPROGDIVRESET (1'b0),
    .CBCC_DATA_SOURCE_SEL ("DECODED"),
    .CDR_SWAP_MODE_EN (1'b0),
    .CHAN_BOND_KEEP_ALIGN ("FALSE"),
    .CHAN_BOND_MAX_SKEW (1),
    .CHAN_BOND_SEQ_1_1 (10'b0000000000),
    .CHAN_BOND_SEQ_1_2 (10'b0000000000),
    .CHAN_BOND_SEQ_1_3 (10'b0000000000),
    .CHAN_BOND_SEQ_1_4 (10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_1 (10'b0000000000),
    .CHAN_BOND_SEQ_2_2 (10'b0000000000),
    .CHAN_BOND_SEQ_2_3 (10'b0000000000),
    .CHAN_BOND_SEQ_2_4 (10'b0000000000),
    .CHAN_BOND_SEQ_2_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_USE ("FALSE"),
    .CHAN_BOND_SEQ_LEN (1),
    .CLK_CORRECT_USE ("FALSE"),
    .CLK_COR_KEEP_IDLE ("FALSE"),
    .CLK_COR_MAX_LAT (12),
    .CLK_COR_MIN_LAT (8),
    .CLK_COR_PRECEDENCE ("TRUE"),
    .CLK_COR_REPEAT_WAIT (0),
    .CLK_COR_SEQ_1_1 (10'b0100000000),
    .CLK_COR_SEQ_1_2 (10'b0100000000),
    .CLK_COR_SEQ_1_3 (10'b0100000000),
    .CLK_COR_SEQ_1_4 (10'b0100000000),
    .CLK_COR_SEQ_1_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_1 (10'b0100000000),
    .CLK_COR_SEQ_2_2 (10'b0100000000),
    .CLK_COR_SEQ_2_3 (10'b0100000000),
    .CLK_COR_SEQ_2_4 (10'b0100000000),
    .CLK_COR_SEQ_2_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_USE ("FALSE"),
    .CLK_COR_SEQ_LEN (1),
    .CPLL_CFG0 (16'h67f8),
    .CPLL_CFG1 (16'ha4ac),
    .CPLL_CFG2 (16'h0007),
    .CPLL_CFG3 (6'h00),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_45 (CPLL_FBDIV_4_5),
    .CPLL_INIT_CFG0 (16'h02b2),
    .CPLL_INIT_CFG1 (8'h00),
    .CPLL_LOCK_CFG (16'h01e8),
    .CPLL_REFCLK_DIV (1),
    .DDI_CTRL (2'b00),
    .DDI_REALIGN_WAIT (15),
    .DEC_MCOMMA_DETECT ("TRUE"),
    .DEC_PCOMMA_DETECT ("TRUE"),
    .DEC_VALID_COMMA_ONLY ("FALSE"),
    .DFE_D_X_REL_POS (1'b0),
    .DFE_VCM_COMP_EN (1'b0),
    .DMONITOR_CFG0 (10'h000),
    .DMONITOR_CFG1 (8'h00),
    .ES_CLK_PHASE_SEL (1'b0),
    .ES_CONTROL (6'b000000),
    .ES_ERRDET_EN ("TRUE"),
    .ES_EYE_SCAN_EN ("TRUE"),
    .ES_HORZ_OFFSET (12'h000),
    .ES_PMA_CFG (10'b0000000000),
    .ES_PRESCALE (5'b00000),
    .ES_QUALIFIER0 (16'h0000),
    .ES_QUALIFIER1 (16'h0000),
    .ES_QUALIFIER2 (16'h0000),
    .ES_QUALIFIER3 (16'h0000),
    .ES_QUALIFIER4 (16'h0000),
    .ES_QUAL_MASK0 (16'h0000),
    .ES_QUAL_MASK1 (16'h0000),
    .ES_QUAL_MASK2 (16'h0000),
    .ES_QUAL_MASK3 (16'h0000),
    .ES_QUAL_MASK4 (16'h0000),
    .ES_SDATA_MASK0 (16'h0000),
    .ES_SDATA_MASK1 (16'h0000),
    .ES_SDATA_MASK2 (16'h0000),
    .ES_SDATA_MASK3 (16'h0000),
    .ES_SDATA_MASK4 (16'h0000),
    .EVODD_PHI_CFG (11'b00000000000),
    .EYE_SCAN_SWAP_EN (1'b0),
    .FTS_DESKEW_SEQ_ENABLE (4'b1111),
    .FTS_LANE_DESKEW_CFG (4'b1111),
    .FTS_LANE_DESKEW_EN ("FALSE"),
    .GEARBOX_MODE (5'b00000),
    .GM_BIAS_SELECT (1'b0),
    .LOCAL_MASTER (1'b1),
    .OOBDIVCTL (2'b00),
    .OOB_PWRUP (1'b0),
    .PCI3_AUTO_REALIGN ("OVR_1K_BLK"),
    .PCI3_PIPE_RX_ELECIDLE (1'b0),
    .PCI3_RX_ASYNC_EBUF_BYPASS (2'b00),
    .PCI3_RX_ELECIDLE_EI2_ENABLE (1'b0),
    .PCI3_RX_ELECIDLE_H2L_COUNT (6'b000000),
    .PCI3_RX_ELECIDLE_H2L_DISABLE (3'b000),
    .PCI3_RX_ELECIDLE_HI_COUNT (6'b000000),
    .PCI3_RX_ELECIDLE_LP4_DISABLE (1'b0),
    .PCI3_RX_FIFO_DISABLE (1'b0),
    .PCIE_BUFG_DIV_CTRL (16'h1000),
    .PCIE_RXPCS_CFG_GEN3 (16'h02a4),
    .PCIE_RXPMA_CFG (16'h000a),
    .PCIE_TXPCS_CFG_GEN3 (16'h24a4),
    .PCIE_TXPMA_CFG (16'h000a),
    .PCS_PCIE_EN ("FALSE"),
    .PCS_RSVD0 (16'b0000000000000000),
    .PCS_RSVD1 (3'b000),
    .PD_TRANS_TIME_FROM_P2 (12'h03c),
    .PD_TRANS_TIME_NONE_P2 (8'h19),
    .PD_TRANS_TIME_TO_P2 (8'h64),
    .PLL_SEL_MODE_GEN12 (2'h3),
    .PLL_SEL_MODE_GEN3 (2'h3),
    .PMA_RSV1 (16'hf000),
    .PROCESS_PAR (3'b010),
    .RATE_SW_USE_DRP (1'b1),
    .RESET_POWERSAVE_DISABLE (1'b0),
    .RXBUFRESET_TIME (5'b00011),
    .RXBUF_ADDR_MODE ("FAST"),
    .RXBUF_EIDLE_HI_CNT (4'b1000),
    .RXBUF_EIDLE_LO_CNT (4'b0000),
    .RXBUF_EN ("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE ("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN ("FALSE"),
    .RXBUF_RESET_ON_EIDLE ("FALSE"),
    .RXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .RXBUF_THRESH_OVFLW (57),
    .RXBUF_THRESH_OVRD ("TRUE"),
    .RXBUF_THRESH_UNDFLW (3),
    .RXCDRFREQRESET_TIME (5'b00001),
    .RXCDRPHRESET_TIME (5'b00001),
    .RXCDR_CFG0 (16'h0000),
    .RXCDR_CFG0_GEN3 (16'h0000),
    .RXCDR_CFG1 (16'h0000),
    .RXCDR_CFG1_GEN3 (16'h0000),
    .RXCDR_CFG2 (16'h0766),
    .RXCDR_CFG2_GEN3 (16'h07e6),
    .RXCDR_CFG3 (16'h0000),
    .RXCDR_CFG3_GEN3 (16'h0000),
    .RXCDR_CFG4 (16'h0000),
    .RXCDR_CFG4_GEN3 (16'h0000),
    .RXCDR_CFG5 (16'h0000),
    .RXCDR_CFG5_GEN3 (16'h0000),
    .RXCDR_FR_RESET_ON_EIDLE (1'b0),
    .RXCDR_HOLD_DURING_EIDLE (1'b0),
    .RXCDR_LOCK_CFG0 (16'h4480),
    .RXCDR_LOCK_CFG1 (16'h5fff),
    .RXCDR_LOCK_CFG2 (16'h77c3),
    .RXCDR_PH_RESET_ON_EIDLE (1'b0),
    .RXCFOK_CFG0 (16'h4000),
    .RXCFOK_CFG1 (16'h0065),
    .RXCFOK_CFG2 (16'h002e),
    .RXDFELPMRESET_TIME (7'b0001111),
    .RXDFELPM_KL_CFG0 (16'h0000),
    .RXDFELPM_KL_CFG1 (16'h0032),
    .RXDFELPM_KL_CFG2 (16'h0000),
    .RXDFE_CFG0 (16'h0a00),
    .RXDFE_CFG1 (16'h0000),
    .RXDFE_GC_CFG0 (16'h0000),
    .RXDFE_GC_CFG1 (16'h7870),
    .RXDFE_GC_CFG2 (16'h0000),
    .RXDFE_H2_CFG0 (16'h0000),
    .RXDFE_H2_CFG1 (16'h0000),
    .RXDFE_H3_CFG0 (16'h4000),
    .RXDFE_H3_CFG1 (16'h0000),
    .RXDFE_H4_CFG0 (16'h2000),
    .RXDFE_H4_CFG1 (16'h0003),
    .RXDFE_H5_CFG0 (16'h2000),
    .RXDFE_H5_CFG1 (16'h0003),
    .RXDFE_H6_CFG0 (16'h2000),
    .RXDFE_H6_CFG1 (16'h0000),
    .RXDFE_H7_CFG0 (16'h2000),
    .RXDFE_H7_CFG1 (16'h0000),
    .RXDFE_H8_CFG0 (16'h2000),
    .RXDFE_H8_CFG1 (16'h0000),
    .RXDFE_H9_CFG0 (16'h2000),
    .RXDFE_H9_CFG1 (16'h0000),
    .RXDFE_HA_CFG0 (16'h2000),
    .RXDFE_HA_CFG1 (16'h0000),
    .RXDFE_HB_CFG0 (16'h2000),
    .RXDFE_HB_CFG1 (16'h0000),
    .RXDFE_HC_CFG0 (16'h0000),
    .RXDFE_HC_CFG1 (16'h0000),
    .RXDFE_HD_CFG0 (16'h0000),
    .RXDFE_HD_CFG1 (16'h0000),
    .RXDFE_HE_CFG0 (16'h0000),
    .RXDFE_HE_CFG1 (16'h0000),
    .RXDFE_HF_CFG0 (16'h0000),
    .RXDFE_HF_CFG1 (16'h0000),
    .RXDFE_OS_CFG0 (16'h8000),
    .RXDFE_OS_CFG1 (16'h0000),
    .RXDFE_UT_CFG0 (16'h8000),
    .RXDFE_UT_CFG1 (16'h0003),
    .RXDFE_VP_CFG0 (16'haa00),
    .RXDFE_VP_CFG1 (16'h0033),
    .RXDLY_CFG (16'h001f),
    .RXDLY_LCFG (16'h0030),
    .RXELECIDLE_CFG ("Sigcfg_4"),
    .RXGBOX_FIFO_INIT_RD_ADDR (4),
    .RXGEARBOX_EN ("FALSE"),
    .RXISCANRESET_TIME (5'b00001),
    .RXLPM_CFG (16'h0000),
    .RXLPM_GC_CFG (16'h1000),
    .RXLPM_KH_CFG0 (16'h0000),
    .RXLPM_KH_CFG1 (16'h0002),
    .RXLPM_OS_CFG0 (16'h8000),
    .RXLPM_OS_CFG1 (16'h0002),
    .RXOOB_CFG (9'b000000110),
    .RXOOB_CLK_CFG ("PMA"),
    .RXOSCALRESET_TIME (5'b00011),
    .RXOUT_DIV (RX_OUT_DIV),
    .RXPCSRESET_TIME (5'b00011),
    .RXPHBEACON_CFG (16'h0000),
    .RXPHDLY_CFG (16'h2020),
    .RXPHSAMP_CFG (16'h2100),
    .RXPHSLIP_CFG (16'h6622),
    .RXPH_MONITOR_SEL (5'b00000),
    .RXPI_CFG0 (2'b01),
    .RXPI_CFG1 (2'b01),
    .RXPI_CFG2 (2'b01),
    .RXPI_CFG3 (2'b01),
    .RXPI_CFG4 (1'b0),
    .RXPI_CFG5 (1'b1),
    .RXPI_CFG6 (3'b011),
    .RXPI_LPM (1'b0),
    .RXPI_VREFSEL (1'b0),
    .RXPMACLK_SEL ("DATA"),
    .RXPMARESET_TIME (5'b00011),
    .RXPRBS_ERR_LOOPBACK (1'b0),
    .RXPRBS_LINKACQ_CNT (15),
    .RXSLIDE_AUTO_WAIT (7),
    .RXSLIDE_MODE ("OFF"),
    .RXSYNC_MULTILANE (1'b1),
    .RXSYNC_OVRD (1'b0),
    .RXSYNC_SKIP_DA (1'b0),
    .RX_AFE_CM_EN (1'b0),
    .RX_BIAS_CFG0 (16'h0ab4),
    .RX_BUFFER_CFG (6'b000000),
    .RX_CAPFF_SARC_ENB (1'b0),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_CLKMUX_EN (1'b1),
    .RX_CLK_SLIP_OVRD (5'b00000),
    .RX_CM_BUF_CFG (4'b1010),
    .RX_CM_BUF_PD (1'b0),
    .RX_CM_SEL (2'b11),
    .RX_CM_TRIM (4'b1010),
    .RX_CTLE3_LPF (8'b00000001),
    .RX_DATA_WIDTH (40),
    .RX_DDI_SEL (6'b000000),
    .RX_DEFER_RESET_BUF_EN ("TRUE"),
    .RX_DFELPM_CFG0 (4'b0110),
    .RX_DFELPM_CFG1 (1'b1),
    .RX_DFELPM_KLKH_AGC_STUP_EN (1'b1),
    .RX_DFE_AGC_CFG0 (2'b10),
    .RX_DFE_AGC_CFG1 (3'b000),
    .RX_DFE_KL_LPM_KH_CFG0 (2'b01),
    .RX_DFE_KL_LPM_KH_CFG1 (3'b000),
    .RX_DFE_KL_LPM_KL_CFG0 (2'b01),
    .RX_DFE_KL_LPM_KL_CFG1 (3'b000),
    .RX_DFE_LPM_HOLD_DURING_EIDLE (1'b0),
    .RX_DISPERR_SEQ_MATCH ("TRUE"),
    .RX_DIVRESET_TIME (5'b00001),
    .RX_EN_HI_LR (1'b1),
    .RX_EYESCAN_VS_CODE (7'b0000000),
    .RX_EYESCAN_VS_NEG_DIR (1'b0),
    .RX_EYESCAN_VS_RANGE (2'b00),
    .RX_EYESCAN_VS_UT_SIGN (1'b0),
    .RX_FABINT_USRCLK_FLOP (1'b0),
    .RX_INT_DATAWIDTH (1),
    .RX_PMA_POWER_SAVE (1'b0),
    .RX_PROGDIV_CFG (0.000000),
    .RX_SAMPLE_PERIOD (3'b111),
    .RX_SIG_VALID_DLY (11),
    .RX_SUM_DFETAPREP_EN (1'b0),
    .RX_SUM_IREF_TUNE (4'b1100),
    .RX_SUM_RES_CTRL (2'b11),
    .RX_SUM_VCMTUNE (4'b0000),
    .RX_SUM_VCM_OVWR (1'b0),
    .RX_SUM_VREF_TUNE (3'b000),
    .RX_TUNE_AFE_OS (2'b10),
    .RX_WIDEMODE_CDR (1'b1),
    .RX_XCLK_SEL ("RXDES"),
    .SAS_MAX_COM (64),
    .SAS_MIN_COM (36),
    .SATA_BURST_SEQ_LEN (4'b1110),
    .SATA_BURST_VAL (3'b100),
    .SATA_CPLL_CFG ("VCO_3000MHZ"),
    .SATA_EIDLE_VAL (3'b100),
    .SATA_MAX_BURST (8),
    .SATA_MAX_INIT (21),
    .SATA_MAX_WAKE (7),
    .SATA_MIN_BURST (4),
    .SATA_MIN_INIT (12),
    .SATA_MIN_WAKE (4),
    .SHOW_REALIGN_COMMA ("TRUE"),
    .SIM_MODE ("FAST"),
    .SIM_RECEIVER_DETECT_PASS ("TRUE"),
    .SIM_RESET_SPEEDUP ("TRUE"),
    .SIM_TX_EIDLE_DRIVE_LEVEL (1'b0),
    .SIM_VERSION (2),
    .TAPDLY_SET_TX (2'h0),
    .TEMPERATUR_PAR (4'b0010),
    .TERM_RCAL_CFG (15'b100001000010000),
    .TERM_RCAL_OVRD (3'b000),
    .TRANS_TIME_RATE (8'h0e),
    .TST_RSV0 (8'h00),
    .TST_RSV1 (8'h00),
    .TXBUF_EN ("TRUE"),
    .TXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .TXDLY_CFG (16'h0009),
    .TXDLY_LCFG (16'h0050),
    .TXDRVBIAS_N (4'b1010),
    .TXDRVBIAS_P (4'b1010),
    .TXFIFO_ADDR_CFG ("LOW"),
    .TXGBOX_FIFO_INIT_RD_ADDR (4),
    .TXGEARBOX_EN ("FALSE"),
    .TXOUT_DIV (TX_OUT_DIV),
    .TXPCSRESET_TIME (5'b00011),
    .TXPHDLY_CFG0 (16'h2020),
    .TXPHDLY_CFG1 (16'h0075),
    .TXPH_CFG (16'h0980),
    .TXPH_MONITOR_SEL (5'b00000),
    .TXPI_CFG0 (2'b01),
    .TXPI_CFG1 (2'b01),
    .TXPI_CFG2 (2'b01),
    .TXPI_CFG3 (1'b0),
    .TXPI_CFG4 (1'b1),
    .TXPI_CFG5 (3'b011),
    .TXPI_GRAY_SEL (1'b0),
    .TXPI_INVSTROBE_SEL (1'b0),
    .TXPI_LPM (1'b0),
    .TXPI_PPMCLK_SEL ("TXUSRCLK2"),
    .TXPI_PPM_CFG (8'b00000000),
    .TXPI_SYNFREQ_PPM (3'b001),
    .TXPI_VREFSEL (1'b0),
    .TXPMARESET_TIME (5'b00011),
    .TXSYNC_MULTILANE (1'b1),
    .TXSYNC_OVRD (1'b0),
    .TXSYNC_SKIP_DA (1'b0),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .TX_CLKMUX_EN (1'b1),
    .TX_DATA_WIDTH (40),
    .TX_DCD_CFG (6'b000010),
    .TX_DCD_EN (1'b0),
    .TX_DEEMPH0 (6'b000000),
    .TX_DEEMPH1 (6'b000000),
    .TX_DIVRESET_TIME (5'b00001),
    .TX_DRIVE_MODE ("DIRECT"),
    .TX_EIDLE_ASSERT_DELAY (3'b100),
    .TX_EIDLE_DEASSERT_DELAY (3'b011),
    .TX_EML_PHI_TUNE (1'b0),
    .TX_FABINT_USRCLK_FLOP (1'b0),
    .TX_IDLE_DATA_ZERO (1'b0),
    .TX_INT_DATAWIDTH (1),
    .TX_LOOPBACK_DRIVE_HIZ ("FALSE"),
    .TX_MAINCURSOR_SEL (1'b0),
    .TX_MARGIN_FULL_0 (7'b1001111),
    .TX_MARGIN_FULL_1 (7'b1001110),
    .TX_MARGIN_FULL_2 (7'b1001100),
    .TX_MARGIN_FULL_3 (7'b1001010),
    .TX_MARGIN_FULL_4 (7'b1001000),
    .TX_MARGIN_LOW_0 (7'b1000110),
    .TX_MARGIN_LOW_1 (7'b1000101),
    .TX_MARGIN_LOW_2 (7'b1000011),
    .TX_MARGIN_LOW_3 (7'b1000010),
    .TX_MARGIN_LOW_4 (7'b1000000),
    .TX_MODE_SEL (3'b000),
    .TX_PMADATA_OPT (1'b0),
    .TX_PMA_POWER_SAVE (1'b0),
    .TX_PROGCLK_SEL ("PREPI"),
    .TX_PROGDIV_CFG (0.000000),
    .TX_QPI_STATUS_EN (1'b0),
    .TX_RXDETECT_CFG (14'h0032),
    .TX_RXDETECT_REF (3'b100),
    .TX_SAMPLE_PERIOD (3'b111),
    .TX_SARC_LPBK_ENB (1'b0),
    .TX_XCLK_SEL ("TXOUT"),
    .USE_PCS_CLK_PHASE_SEL (1'b0),
    .WB_MODE (2'b00))
  i_gthe3_channel (
    .BUFGTCE (),
    .BUFGTCEMASK (),
    .BUFGTDIV (),
    .BUFGTRESET (),
    .BUFGTRSTMASK (),
    .CFGRESET (1'h0),
    .CLKRSVD0 (1'h0),
    .CLKRSVD1 (1'h0),
    .CPLLFBCLKLOST (),
    .CPLLLOCK (cpll_locked_s),
    .CPLLLOCKDETCLK (up_clk),
    .CPLLLOCKEN (1'h1),
    .CPLLPD (1'h0),
    .CPLLREFCLKLOST (),
    .CPLLREFCLKSEL (3'h1),
    .CPLLRESET (up_cpll_rst),
    .DMONFIFORESET (1'h0),
    .DMONITORCLK (1'h0),
    .DMONITOROUT (),
    .DRPADDR (up_addr_int[8:0]),
    .DRPCLK (up_clk),
    .DRPDI (up_wdata_int),
    .DRPDO (up_rdata_s),
    .DRPEN (up_enb_int),
    .DRPRDY (up_ready_s),
    .DRPWE (up_wr_int),
    .EVODDPHICALDONE (1'h0),
    .EVODDPHICALSTART (1'h0),
    .EVODDPHIDRDEN (1'h0),
    .EVODDPHIDWREN (1'h0),
    .EVODDPHIXRDEN (1'h0),
    .EVODDPHIXWREN (1'h0),
    .EYESCANDATAERROR (),
    .EYESCANMODE (1'h0),
    .EYESCANRESET (1'h0),
    .EYESCANTRIGGER (1'h0),
    .GTGREFCLK (1'h0),
    .GTHRXN (rx_n),
    .GTHRXP (rx_p),
    .GTHTXN (tx_n),
    .GTHTXP (tx_p),
    .GTNORTHREFCLK0 (1'h0),
    .GTNORTHREFCLK1 (1'h0),
    .GTPOWERGOOD (),
    .GTREFCLK0 (cpll_ref_clk),
    .GTREFCLK1 (1'h0),
    .GTREFCLKMONITOR (),
    .GTRESETSEL (1'h0),
    .GTRSVD (16'h0),
    .GTRXRESET (up_rx_rst),
    .GTSOUTHREFCLK0 (1'h0),
    .GTSOUTHREFCLK1 (1'h0),
    .GTTXRESET (up_tx_rst),
    .LOOPBACK (3'h0),
    .LPBKRXTXSEREN (1'h0),
    .LPBKTXRXSEREN (1'h0),
    .PCIEEQRXEQADAPTDONE (1'h0),
    .PCIERATEGEN3 (),
    .PCIERATEIDLE (),
    .PCIERATEQPLLPD (),
    .PCIERATEQPLLRESET (),
    .PCIERSTIDLE (1'h0),
    .PCIERSTTXSYNCSTART (1'h0),
    .PCIESYNCTXSYNCDONE (),
    .PCIEUSERGEN3RDY (),
    .PCIEUSERPHYSTATUSRST (),
    .PCIEUSERRATEDONE (1'h0),
    .PCIEUSERRATESTART (),
    .PCSRSVDIN (16'h0),
    .PCSRSVDIN2 (5'h0),
    .PCSRSVDOUT (),
    .PHYSTATUS (),
    .PINRSRVDAS (),
    .PMARSVDIN (5'h0),
    .QPLL0CLK (qpll2ch_clk),
    .QPLL0REFCLK (qpll2ch_ref_clk),
    .QPLL1CLK (1'h0),
    .QPLL1REFCLK (1'h0),
    .RESETEXCEPTION (),
    .RESETOVRD (1'h0),
    .RSTCLKENTX (1'h0),
    .RX8B10BEN (1'h1),
    .RXBUFRESET (1'h0),
    .RXBUFSTATUS (),
    .RXBYTEISALIGNED (),
    .RXBYTEREALIGN (),
    .RXCDRFREQRESET (1'h0),
    .RXCDRHOLD (1'h0),
    .RXCDRLOCK (),
    .RXCDROVRDEN (1'h0),
    .RXCDRPHDONE (),
    .RXCDRRESET (1'h0),
    .RXCDRRESETRSV (1'h0),
    .RXCHANBONDSEQ (),
    .RXCHANISALIGNED (),
    .RXCHANREALIGN (),
    .RXCHBONDEN (1'h0),
    .RXCHBONDI (5'h0),
    .RXCHBONDLEVEL (3'h0),
    .RXCHBONDMASTER (1'h0),
    .RXCHBONDO (),
    .RXCHBONDSLAVE (1'h0),
    .RXCLKCORCNT (),
    .RXCOMINITDET (),
    .RXCOMMADET (),
    .RXCOMMADETEN (1'h1),
    .RXCOMSASDET (),
    .RXCOMWAKEDET (),
    .RXCTRL0 ({rx_charisk_open_s, rx_charisk}),
    .RXCTRL1 ({rx_disperr_open_s, rx_disperr}),
    .RXCTRL2 (),
    .RXCTRL3 ({rx_notintable_open_s, rx_notintable}),
    .RXDATA ({rx_data_open_s, rx_data}),
    .RXDATAEXTENDRSVD (),
    .RXDATAVALID (),
    .RXDFEAGCCTRL (2'h1),
    .RXDFEAGCHOLD (1'h0),
    .RXDFEAGCOVRDEN (1'h0),
    .RXDFELFHOLD (1'h0),
    .RXDFELFOVRDEN (1'h0),
    .RXDFELPMRESET (1'h0),
    .RXDFETAP10HOLD (1'h0),
    .RXDFETAP10OVRDEN (1'h0),
    .RXDFETAP11HOLD (1'h0),
    .RXDFETAP11OVRDEN (1'h0),
    .RXDFETAP12HOLD (1'h0),
    .RXDFETAP12OVRDEN (1'h0),
    .RXDFETAP13HOLD (1'h0),
    .RXDFETAP13OVRDEN (1'h0),
    .RXDFETAP14HOLD (1'h0),
    .RXDFETAP14OVRDEN (1'h0),
    .RXDFETAP15HOLD (1'h0),
    .RXDFETAP15OVRDEN (1'h0),
    .RXDFETAP2HOLD (1'h0),
    .RXDFETAP2OVRDEN (1'h0),
    .RXDFETAP3HOLD (1'h0),
    .RXDFETAP3OVRDEN (1'h0),
    .RXDFETAP4HOLD (1'h0),
    .RXDFETAP4OVRDEN (1'h0),
    .RXDFETAP5HOLD (1'h0),
    .RXDFETAP5OVRDEN (1'h0),
    .RXDFETAP6HOLD (1'h0),
    .RXDFETAP6OVRDEN (1'h0),
    .RXDFETAP7HOLD (1'h0),
    .RXDFETAP7OVRDEN (1'h0),
    .RXDFETAP8HOLD (1'h0),
    .RXDFETAP8OVRDEN (1'h0),
    .RXDFETAP9HOLD (1'h0),
    .RXDFETAP9OVRDEN (1'h0),
    .RXDFEUTHOLD (1'h0),
    .RXDFEUTOVRDEN (1'h0),
    .RXDFEVPHOLD (1'h0),
    .RXDFEVPOVRDEN (1'h0),
    .RXDFEVSEN (1'h0),
    .RXDFEXYDEN (1'h1),
    .RXDLYBYPASS (1'h1),
    .RXDLYEN (1'h0),
    .RXDLYOVRDEN (1'h0),
    .RXDLYSRESET (1'h0),
    .RXDLYSRESETDONE (),
    .RXELECIDLE (),
    .RXELECIDLEMODE (2'h3),
    .RXGEARBOXSLIP (1'h0),
    .RXHEADER (),
    .RXHEADERVALID (),
    .RXLATCLK (1'h0),
    .RXLPMEN (up_rx_lpm_dfe_n),
    .RXLPMGCHOLD (1'h0),
    .RXLPMGCOVRDEN (1'h0),
    .RXLPMHFHOLD (1'h0),
    .RXLPMHFOVRDEN (1'h0),
    .RXLPMLFHOLD (1'h0),
    .RXLPMLFKLOVRDEN (1'h0),
    .RXLPMOSHOLD (1'h0),
    .RXLPMOSOVRDEN (1'h0),
    .RXMCOMMAALIGNEN (rx_calign),
    .RXMONITOROUT (),
    .RXMONITORSEL (2'h0),
    .RXOOBRESET (1'h0),
    .RXOSCALRESET (1'h0),
    .RXOSHOLD (1'h0),
    .RXOSINTCFG (4'hd),
    .RXOSINTDONE (),
    .RXOSINTEN (1'h1),
    .RXOSINTHOLD (1'h0),
    .RXOSINTOVRDEN (1'h0),
    .RXOSINTSTARTED (),
    .RXOSINTSTROBE (1'h0),
    .RXOSINTSTROBEDONE (),
    .RXOSINTSTROBESTARTED (),
    .RXOSINTTESTOVRDEN (1'h0),
    .RXOSOVRDEN (1'h0),
    .RXOUTCLK (rx_out_clk_s),
    .RXOUTCLKFABRIC (),
    .RXOUTCLKPCS (),
    .RXOUTCLKSEL (up_rx_out_clk_sel),
    .RXPCOMMAALIGNEN (rx_calign),
    .RXPCSRESET (1'h0),
    .RXPD (2'h0),
    .RXPHALIGN (1'h0),
    .RXPHALIGNDONE (),
    .RXPHALIGNEN (1'h0),
    .RXPHALIGNERR (),
    .RXPHDLYPD (1'h1),
    .RXPHDLYRESET (1'h0),
    .RXPHOVRDEN (1'h0),
    .RXPLLCLKSEL (rx_pll_clk_sel_s),
    .RXPMARESET (1'h0),
    .RXPMARESETDONE (),
    .RXPOLARITY (1'h0),
    .RXPRBSCNTRESET (1'h0),
    .RXPRBSERR (),
    .RXPRBSLOCKED (),
    .RXPRBSSEL (4'h0),
    .RXPRGDIVRESETDONE (),
    .RXPROGDIVRESET (1'h0),
    .RXQPIEN (1'h0),
    .RXQPISENN (),
    .RXQPISENP (),
    .RXRATE (rx_rate_m2),
    .RXRATEDONE (),
    .RXRATEMODE (1'h0),
    .RXRECCLKOUT (),
    .RXRESETDONE (rx_rst_done_s),
    .RXSLIDE (1'h0),
    .RXSLIDERDY (),
    .RXSLIPDONE (),
    .RXSLIPOUTCLK (1'h0),
    .RXSLIPOUTCLKRDY (),
    .RXSLIPPMA (1'h0),
    .RXSLIPPMARDY (),
    .RXSTARTOFSEQ (),
    .RXSTATUS (),
    .RXSYNCALLIN (1'h0),
    .RXSYNCDONE (),
    .RXSYNCIN (1'h0),
    .RXSYNCMODE (1'h0),
    .RXSYNCOUT (),
    .RXSYSCLKSEL (rx_sys_clk_sel_s),
    .RXUSERRDY (up_rx_user_ready),
    .RXUSRCLK (rx_clk),
    .RXUSRCLK2 (rx_clk),
    .RXVALID (),
    .SIGVALIDCLK (1'h0),
    .TSTIN (20'h0),
    .TX8B10BBYPASS (8'h0),
    .TX8B10BEN (1'h1),
    .TXBUFDIFFCTRL (3'h0),
    .TXBUFSTATUS (),
    .TXCOMFINISH (),
    .TXCOMINIT (1'h0),
    .TXCOMSAS (1'h0),
    .TXCOMWAKE (1'h0),
    .TXCTRL0 (16'h0),
    .TXCTRL1 (16'h0),
    .TXCTRL2 ({4'd0, tx_charisk}),
    .TXDATA ({96'd0, tx_data}),
    .TXDATAEXTENDRSVD (8'h0),
    .TXDEEMPH (1'h0),
    .TXDETECTRX (1'h0),
    .TXDIFFCTRL (4'h8),
    .TXDIFFPD (1'h0),
    .TXDLYBYPASS (1'h1),
    .TXDLYEN (1'h0),
    .TXDLYHOLD (1'h0),
    .TXDLYOVRDEN (1'h0),
    .TXDLYSRESET (1'h0),
    .TXDLYSRESETDONE (),
    .TXDLYUPDOWN (1'h0),
    .TXELECIDLE (1'h0),
    .TXHEADER (6'h0),
    .TXINHIBIT (1'h0),
    .TXLATCLK (1'h0),
    .TXMAINCURSOR (7'h40),
    .TXMARGIN (3'h0),
    .TXOUTCLK (tx_out_clk_s),
    .TXOUTCLKFABRIC (),
    .TXOUTCLKPCS (),
    .TXOUTCLKSEL (up_tx_out_clk_sel),
    .TXPCSRESET (1'h0),
    .TXPD (2'h0),
    .TXPDELECIDLEMODE (1'h0),
    .TXPHALIGN (1'h0),
    .TXPHALIGNDONE (),
    .TXPHALIGNEN (1'h0),
    .TXPHDLYPD (1'h1),
    .TXPHDLYRESET (1'h0),
    .TXPHDLYTSTCLK (1'h0),
    .TXPHINIT (1'h0),
    .TXPHINITDONE (),
    .TXPHOVRDEN (1'h0),
    .TXPIPPMEN (1'h0),
    .TXPIPPMOVRDEN (1'h0),
    .TXPIPPMPD (1'h0),
    .TXPIPPMSEL (1'h0),
    .TXPIPPMSTEPSIZE (5'h0),
    .TXPISOPD (1'h0),
    .TXPLLCLKSEL (tx_pll_clk_sel_s),
    .TXPMARESET (1'h0),
    .TXPMARESETDONE (),
    .TXPOLARITY (1'h0),
    .TXPOSTCURSOR (5'h0),
    .TXPOSTCURSORINV (1'h0),
    .TXPRBSFORCEERR (1'h0),
    .TXPRBSSEL (4'h0),
    .TXPRECURSOR (5'h0),
    .TXPRECURSORINV (1'h0),
    .TXPRGDIVRESETDONE (),
    .TXPROGDIVRESET (up_tx_rst),
    .TXQPIBIASEN (1'h0),
    .TXQPISENN (),
    .TXQPISENP (),
    .TXQPISTRONGPDOWN (1'h0),
    .TXQPIWEAKPUP (1'h0),
    .TXRATE (tx_rate_m2),
    .TXRATEDONE (),
    .TXRATEMODE (1'h0),
    .TXRESETDONE (tx_rst_done_s),
    .TXSEQUENCE (7'h0),
    .TXSWING (1'h0),
    .TXSYNCALLIN (1'h0),
    .TXSYNCDONE (),
    .TXSYNCIN (1'h0),
    .TXSYNCMODE (1'h0),
    .TXSYNCOUT (),
    .TXSYSCLKSEL (tx_sys_clk_sel_s),
    .TXUSERRDY (up_tx_user_ready),
    .TXUSRCLK (tx_clk),
    .TXUSRCLK2 (tx_clk));
  end
  endgenerate

  generate
  if (XCVR_TYPE == 2) begin
  BUFG_GT i_rx_bufg (
    .CE (1'b1),
    .CEMASK (1'b0),
    .CLR (1'b0),
    .CLRMASK (1'b0),
    .DIV (3'd0),
    .I (rx_out_clk_s),
    .O (rx_out_clk));

  BUFG_GT i_tx_bufg (
    .CE (1'b1),
    .CEMASK (1'b0),
    .CLR (1'b0),
    .CLRMASK (1'b0),
    .DIV (3'd0),
    .I (tx_out_clk_s),
    .O (tx_out_clk));
  end
  endgenerate

  generate
  if (XCVR_TYPE == 2) begin
  assign rx_sys_clk_sel_s = (up_rx_sys_clk_sel == 2'd3) ? 2'b10 : 2'b00;
  assign tx_sys_clk_sel_s = (up_tx_sys_clk_sel == 2'd3) ? 2'b10 : 2'b00;
  assign rx_pll_clk_sel_s = up_rx_sys_clk_sel;
  assign tx_pll_clk_sel_s = up_tx_sys_clk_sel;
  end
  endgenerate

  generate
  if (XCVR_TYPE == 2) begin
  GTHE4_CHANNEL #(
    .ACJTAG_DEBUG_MODE (1'b0),
    .ACJTAG_MODE (1'b0),
    .ACJTAG_RESET (1'b0),
    .ADAPT_CFG0 (16'h1000),
    .ADAPT_CFG1 (16'hc800),
    .ADAPT_CFG2 (16'h0000),
    .ALIGN_COMMA_DOUBLE ("FALSE"),
    .ALIGN_COMMA_ENABLE (10'b1111111111),
    .ALIGN_COMMA_WORD (1'h1),
    .ALIGN_MCOMMA_DET ("TRUE"),
    .ALIGN_MCOMMA_VALUE (10'b1010000011),
    .ALIGN_PCOMMA_DET ("TRUE"),
    .ALIGN_PCOMMA_VALUE (10'b0101111100),
    .A_RXOSCALRESET (1'b0),
    .A_RXPROGDIVRESET (1'b0),
    .A_RXTERMINATION (1'b1),
    .A_TXDIFFCTRL (5'b01100),
    .A_TXPROGDIVRESET (1'b0),
    .CAPBYPASS_FORCE (1'b0),
    .CBCC_DATA_SOURCE_SEL ("DECODED"),
    .CDR_SWAP_MODE_EN (1'b0),
    .CFOK_PWRSVE_EN (1'b1),
    .CHAN_BOND_KEEP_ALIGN ("FALSE"),
    .CHAN_BOND_MAX_SKEW (1'h1),
    .CHAN_BOND_SEQ_1_1 (10'b0000000000),
    .CHAN_BOND_SEQ_1_2 (10'b0000000000),
    .CHAN_BOND_SEQ_1_3 (10'b0000000000),
    .CHAN_BOND_SEQ_1_4 (10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_1 (10'b0000000000),
    .CHAN_BOND_SEQ_2_2 (10'b0000000000),
    .CHAN_BOND_SEQ_2_3 (10'b0000000000),
    .CHAN_BOND_SEQ_2_4 (10'b0000000000),
    .CHAN_BOND_SEQ_2_ENABLE (4'b1111),
    .CHAN_BOND_SEQ_2_USE ("FALSE"),
    .CHAN_BOND_SEQ_LEN (1'h1),
    .CH_HSPMUX (16'h2424),
    .CKCAL1_CFG_0 (16'b1100000011000000),
    .CKCAL1_CFG_1 (16'b0101000011000000),
    .CKCAL1_CFG_2 (16'b0000000000001010),
    .CKCAL1_CFG_3 (16'b0000000000000000),
    .CKCAL2_CFG_0 (16'b1100000011000000),
    .CKCAL2_CFG_1 (16'b1000000011000000),
    .CKCAL2_CFG_2 (16'b0000000000000000),
    .CKCAL2_CFG_3 (16'b0000000000000000),
    .CKCAL2_CFG_4 (16'b0000000000000000),
    .CKCAL_RSVD0 (16'h0080),
    .CKCAL_RSVD1 (16'h0400),
    .CLK_CORRECT_USE ("FALSE"),
    .CLK_COR_KEEP_IDLE ("FALSE"),
    .CLK_COR_MAX_LAT (12),
    .CLK_COR_MIN_LAT (8),
    .CLK_COR_PRECEDENCE ("TRUE"),
    .CLK_COR_REPEAT_WAIT (1'h0),
    .CLK_COR_SEQ_1_1 (10'b0100000000),
    .CLK_COR_SEQ_1_2 (10'b0100000000),
    .CLK_COR_SEQ_1_3 (10'b0100000000),
    .CLK_COR_SEQ_1_4 (10'b0100000000),
    .CLK_COR_SEQ_1_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_1 (10'b0100000000),
    .CLK_COR_SEQ_2_2 (10'b0100000000),
    .CLK_COR_SEQ_2_3 (10'b0100000000),
    .CLK_COR_SEQ_2_4 (10'b0100000000),
    .CLK_COR_SEQ_2_ENABLE (4'b1111),
    .CLK_COR_SEQ_2_USE ("FALSE"),
    .CLK_COR_SEQ_LEN (1'h1),
    .CPLL_CFG0 (16'h01fa),
    .CPLL_CFG1 (16'h0023),
    .CPLL_CFG2 (16'h0002),
    .CPLL_CFG3 (16'h0000),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_45 (5),
    .CPLL_INIT_CFG0 (16'h02b2),
    .CPLL_LOCK_CFG (16'h01e8),
    .CPLL_REFCLK_DIV (1'h1),
    .CTLE3_OCAP_EXT_CTRL (3'b000),
    .CTLE3_OCAP_EXT_EN (1'b0),
    .DDI_CTRL (2'b00),
    .DDI_REALIGN_WAIT (15),
    .DEC_MCOMMA_DETECT ("TRUE"),
    .DEC_PCOMMA_DETECT ("TRUE"),
    .DEC_VALID_COMMA_ONLY ("FALSE"),
    .DELAY_ELEC (1'b0),
    .DMONITOR_CFG0 (10'h000),
    .DMONITOR_CFG1 (8'h00),
    .ES_CLK_PHASE_SEL (1'b0),
    .ES_CONTROL (6'b000000),
    .ES_ERRDET_EN ("TRUE"),
    .ES_EYE_SCAN_EN ("TRUE"),
    .ES_HORZ_OFFSET (12'h000),
    .ES_PRESCALE (5'b00000),
    .ES_QUALIFIER0 (16'h0000),
    .ES_QUALIFIER1 (16'h0000),
    .ES_QUALIFIER2 (16'h0000),
    .ES_QUALIFIER3 (16'h0000),
    .ES_QUALIFIER4 (16'h0000),
    .ES_QUALIFIER5 (16'h0000),
    .ES_QUALIFIER6 (16'h0000),
    .ES_QUALIFIER7 (16'h0000),
    .ES_QUALIFIER8 (16'h0000),
    .ES_QUALIFIER9 (16'h0000),
    .ES_QUAL_MASK0 (16'h0000),
    .ES_QUAL_MASK1 (16'h0000),
    .ES_QUAL_MASK2 (16'h0000),
    .ES_QUAL_MASK3 (16'h0000),
    .ES_QUAL_MASK4 (16'h0000),
    .ES_QUAL_MASK5 (16'h0000),
    .ES_QUAL_MASK6 (16'h0000),
    .ES_QUAL_MASK7 (16'h0000),
    .ES_QUAL_MASK8 (16'h0000),
    .ES_QUAL_MASK9 (16'h0000),
    .ES_SDATA_MASK0 (16'h0000),
    .ES_SDATA_MASK1 (16'h0000),
    .ES_SDATA_MASK2 (16'h0000),
    .ES_SDATA_MASK3 (16'h0000),
    .ES_SDATA_MASK4 (16'h0000),
    .ES_SDATA_MASK5 (16'h0000),
    .ES_SDATA_MASK6 (16'h0000),
    .ES_SDATA_MASK7 (16'h0000),
    .ES_SDATA_MASK8 (16'h0000),
    .ES_SDATA_MASK9 (16'h0000),
    .EYE_SCAN_SWAP_EN (1'b0),
    .FTS_DESKEW_SEQ_ENABLE (4'b1111),
    .FTS_LANE_DESKEW_CFG (4'b1111),
    .FTS_LANE_DESKEW_EN ("FALSE"),
    .GEARBOX_MODE (5'b00000),
    .ISCAN_CK_PH_SEL2 (1'b0),
    .LOCAL_MASTER (1'b1),
    .LPBK_BIAS_CTRL (3'b100),
    .LPBK_EN_RCAL_B (1'b0),
    .LPBK_EXT_RCAL (4'b1000),
    .LPBK_IND_CTRL0 (3'b000),
    .LPBK_IND_CTRL1 (3'b000),
    .LPBK_IND_CTRL2 (3'b000),
    .LPBK_RG_CTRL (4'b1110),
    .OOBDIVCTL (2'b00),
    .OOB_PWRUP (1'b0),
    .PCI3_AUTO_REALIGN ("OVR_1K_BLK"),
    .PCI3_PIPE_RX_ELECIDLE (1'b0),
    .PCI3_RX_ASYNC_EBUF_BYPASS (2'b00),
    .PCI3_RX_ELECIDLE_EI2_ENABLE (1'b0),
    .PCI3_RX_ELECIDLE_H2L_COUNT (6'b000000),
    .PCI3_RX_ELECIDLE_H2L_DISABLE (3'b000),
    .PCI3_RX_ELECIDLE_HI_COUNT (6'b000000),
    .PCI3_RX_ELECIDLE_LP4_DISABLE (1'b0),
    .PCI3_RX_FIFO_DISABLE (1'b0),
    .PCIE3_CLK_COR_EMPTY_THRSH (5'b00000),
    .PCIE3_CLK_COR_FULL_THRSH (6'b010000),
    .PCIE3_CLK_COR_MAX_LAT (5'b00100),
    .PCIE3_CLK_COR_MIN_LAT (5'b00000),
    .PCIE3_CLK_COR_THRSH_TIMER (6'b001000),
    .PCIE_BUFG_DIV_CTRL (16'h3500),
    .PCIE_PLL_SEL_MODE_GEN12 (2'h2),
    .PCIE_PLL_SEL_MODE_GEN3 (2'h2),
    .PCIE_PLL_SEL_MODE_GEN4 (2'h2),
    .PCIE_RXPCS_CFG_GEN3 (16'h0aa5),
    .PCIE_RXPMA_CFG (16'h280a),
    .PCIE_TXPCS_CFG_GEN3 (16'h24a4),
    .PCIE_TXPMA_CFG (16'h280a),
    .PCS_PCIE_EN ("FALSE"),
    .PCS_RSVD0 (16'b0000000000000000),
    .PD_TRANS_TIME_FROM_P2 (12'h03c),
    .PD_TRANS_TIME_NONE_P2 (8'h19),
    .PD_TRANS_TIME_TO_P2 (8'h64),
    .PREIQ_FREQ_BST (1'h0),
    .PROCESS_PAR (3'b010),
    .RATE_SW_USE_DRP (1'b1),
    .RCLK_SIPO_DLY_ENB (1'b0),
    .RCLK_SIPO_INV_EN (1'b0),
    .RESET_POWERSAVE_DISABLE (1'b0),
    .RTX_BUF_CML_CTRL (3'b010),
    .RTX_BUF_TERM_CTRL (2'b00),
    .RXBUFRESET_TIME (5'b00011),
    .RXBUF_ADDR_MODE ("FAST"),
    .RXBUF_EIDLE_HI_CNT (4'b1000),
    .RXBUF_EIDLE_LO_CNT (4'b0000),
    .RXBUF_EN ("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE ("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN ("FALSE"),
    .RXBUF_RESET_ON_EIDLE ("FALSE"),
    .RXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .RXBUF_THRESH_OVFLW (57),
    .RXBUF_THRESH_OVRD ("TRUE"),
    .RXBUF_THRESH_UNDFLW (3),
    .RXCDRFREQRESET_TIME (5'b00001),
    .RXCDRPHRESET_TIME (5'b00001),
    .RXCDR_CFG0 (16'h0002),
    .RXCDR_CFG0_GEN3 (16'h0003),
    .RXCDR_CFG1 (16'h0000),
    .RXCDR_CFG1_GEN3 (16'h0000),
    .RXCDR_CFG2 (16'h0265),
    .RXCDR_CFG2_GEN3 (16'h0265),
    .RXCDR_CFG2_GEN4 (16'h00b4),
    .RXCDR_CFG3 (16'h0012),
    .RXCDR_CFG3_GEN3 (16'h0012),
    .RXCDR_CFG3_GEN4 (16'h0024),
    .RXCDR_CFG4 (16'h5cf6),
    .RXCDR_CFG4_GEN3 (16'h5cf6),
    .RXCDR_CFG5 (16'hb46b),
    .RXCDR_CFG5_GEN3 (16'h146b),
    .RXCDR_FR_RESET_ON_EIDLE (1'b0),
    .RXCDR_HOLD_DURING_EIDLE (1'b0),
    .RXCDR_LOCK_CFG0 (16'h2201),
    .RXCDR_LOCK_CFG1 (16'h9fff),
    .RXCDR_LOCK_CFG2 (16'h77c3),
    .RXCDR_LOCK_CFG3 (16'h0001),
    .RXCDR_LOCK_CFG4 (16'h0000),
    .RXCDR_PH_RESET_ON_EIDLE (1'b0),
    .RXCFOK_CFG0 (16'h0000),
    .RXCFOK_CFG1 (16'h8015),
    .RXCFOK_CFG2 (16'h02ae),
    .RXCKCAL1_IQ_LOOP_RST_CFG (16'h0004),
    .RXCKCAL1_I_LOOP_RST_CFG (16'h0004),
    .RXCKCAL1_Q_LOOP_RST_CFG (16'h0004),
    .RXCKCAL2_DX_LOOP_RST_CFG (16'h0004),
    .RXCKCAL2_D_LOOP_RST_CFG (16'h0004),
    .RXCKCAL2_S_LOOP_RST_CFG (16'h0004),
    .RXCKCAL2_X_LOOP_RST_CFG (16'h0004),
    .RXDFELPMRESET_TIME (7'b0001111),
    .RXDFELPM_KL_CFG0 (16'h0000),
    .RXDFELPM_KL_CFG1 (16'ha0e2),
    .RXDFELPM_KL_CFG2 (16'h0100),
    .RXDFE_CFG0 (16'h0a00),
    .RXDFE_CFG1 (16'h0280),
    .RXDFE_GC_CFG0 (16'h0000),
    .RXDFE_GC_CFG1 (16'h8000),
    .RXDFE_GC_CFG2 (16'hffe0),
    .RXDFE_H2_CFG0 (16'h0000),
    .RXDFE_H2_CFG1 (16'h0002),
    .RXDFE_H3_CFG0 (16'h0000),
    .RXDFE_H3_CFG1 (16'h8002),
    .RXDFE_H4_CFG0 (16'h0000),
    .RXDFE_H4_CFG1 (16'h8002),
    .RXDFE_H5_CFG0 (16'h0000),
    .RXDFE_H5_CFG1 (16'h8002),
    .RXDFE_H6_CFG0 (16'h0000),
    .RXDFE_H6_CFG1 (16'h8002),
    .RXDFE_H7_CFG0 (16'h0000),
    .RXDFE_H7_CFG1 (16'h8002),
    .RXDFE_H8_CFG0 (16'h0000),
    .RXDFE_H8_CFG1 (16'h8002),
    .RXDFE_H9_CFG0 (16'h0000),
    .RXDFE_H9_CFG1 (16'h8002),
    .RXDFE_HA_CFG0 (16'h0000),
    .RXDFE_HA_CFG1 (16'h8002),
    .RXDFE_HB_CFG0 (16'h0000),
    .RXDFE_HB_CFG1 (16'h8002),
    .RXDFE_HC_CFG0 (16'h0000),
    .RXDFE_HC_CFG1 (16'h8002),
    .RXDFE_HD_CFG0 (16'h0000),
    .RXDFE_HD_CFG1 (16'h8002),
    .RXDFE_HE_CFG0 (16'h0000),
    .RXDFE_HE_CFG1 (16'h8002),
    .RXDFE_HF_CFG0 (16'h0000),
    .RXDFE_HF_CFG1 (16'h8002),
    .RXDFE_KH_CFG0 (16'h0000),
    .RXDFE_KH_CFG1 (16'h8000),
    .RXDFE_KH_CFG2 (16'h2613),
    .RXDFE_KH_CFG3 (16'h411c),
    .RXDFE_OS_CFG0 (16'h0000),
    .RXDFE_OS_CFG1 (16'h8002),
    .RXDFE_PWR_SAVING (1'b1),
    .RXDFE_UT_CFG0 (16'h0000),
    .RXDFE_UT_CFG1 (16'h0003),
    .RXDFE_UT_CFG2 (16'h0000),
    .RXDFE_VP_CFG0 (16'h0000),
    .RXDFE_VP_CFG1 (16'h8033),
    .RXDLY_CFG (16'h0010),
    .RXDLY_LCFG (16'h0030),
    .RXELECIDLE_CFG ("SIGCFG_4"),
    .RXGBOX_FIFO_INIT_RD_ADDR (4),
    .RXGEARBOX_EN ("FALSE"),
    .RXISCANRESET_TIME (5'b00001),
    .RXLPM_CFG (16'h0000),
    .RXLPM_GC_CFG (16'h8000),
    .RXLPM_KH_CFG0 (16'h0000),
    .RXLPM_KH_CFG1 (16'h0002),
    .RXLPM_OS_CFG0 (16'h0000),
    .RXLPM_OS_CFG1 (16'h8002),
    .RXOOB_CFG (9'b000000110),
    .RXOOB_CLK_CFG ("PMA"),
    .RXOSCALRESET_TIME (5'b00011),
    .RXOUT_DIV (RX_OUT_DIV),
    .RXPCSRESET_TIME (5'b00011),
    .RXPHBEACON_CFG (16'h0000),
    .RXPHDLY_CFG (16'h2070),
    .RXPHSAMP_CFG (16'h2100),
    .RXPHSLIP_CFG (16'h9933),
    .RXPH_MONITOR_SEL (5'b00000),
    .RXPI_AUTO_BW_SEL_BYPASS (1'b0),
    .RXPI_CFG0 (16'h0002),
    .RXPI_CFG1 (16'b0000000000010101),
    .RXPI_LPM (1'b0),
    .RXPI_SEL_LC (2'b00),
    .RXPI_STARTCODE (2'b00),
    .RXPI_VREFSEL (1'b0),
    .RXPMACLK_SEL ("DATA"),
    .RXPMARESET_TIME (5'b00011),
    .RXPRBS_ERR_LOOPBACK (1'b0),
    .RXPRBS_LINKACQ_CNT (15),
    .RXREFCLKDIV2_SEL (1'b0),
    .RXSLIDE_AUTO_WAIT (7),
    .RXSLIDE_MODE ("OFF"),
    .RXSYNC_MULTILANE (1'b1),
    .RXSYNC_OVRD (1'b0),
    .RXSYNC_SKIP_DA (1'b0),
    .RX_AFE_CM_EN (1'b0),
    .RX_BIAS_CFG0 (16'h1554),
    .RX_BUFFER_CFG (6'b000000),
    .RX_CAPFF_SARC_ENB (1'b0),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_CLKMUX_EN (1'b1),
    .RX_CLK_SLIP_OVRD (5'b00000),
    .RX_CM_BUF_CFG (4'b1010),
    .RX_CM_BUF_PD (1'b0),
    .RX_CM_SEL (3),
    .RX_CM_TRIM (10),
    .RX_CTLE3_LPF (8'b11111111),
    .RX_DATA_WIDTH (40),
    .RX_DDI_SEL (6'b000000),
    .RX_DEFER_RESET_BUF_EN ("TRUE"),
    .RX_DEGEN_CTRL (3'b011),
    .RX_DFELPM_CFG0 (6),
    .RX_DFELPM_CFG1 (1'b1),
    .RX_DFELPM_KLKH_AGC_STUP_EN (1'b1),
    .RX_DFE_AGC_CFG0 (2'b10),
    .RX_DFE_AGC_CFG1 (4),
    .RX_DFE_KL_LPM_KH_CFG0 (1'h1),
    .RX_DFE_KL_LPM_KH_CFG1 (4),
    .RX_DFE_KL_LPM_KL_CFG0 (2'b01),
    .RX_DFE_KL_LPM_KL_CFG1 (4),
    .RX_DFE_LPM_HOLD_DURING_EIDLE (1'b0),
    .RX_DISPERR_SEQ_MATCH ("TRUE"),
    .RX_DIV2_MODE_B (1'b0),
    .RX_DIVRESET_TIME (5'b00001),
    .RX_EN_CTLE_RCAL_B (1'b0),
    .RX_EN_HI_LR (1'b1),
    .RX_EXT_RL_CTRL (9'b000000000),
    .RX_EYESCAN_VS_CODE (7'b0000000),
    .RX_EYESCAN_VS_NEG_DIR (1'b0),
    .RX_EYESCAN_VS_RANGE (2'b00),
    .RX_EYESCAN_VS_UT_SIGN (1'b0),
    .RX_FABINT_USRCLK_FLOP (1'b0),
    .RX_INT_DATAWIDTH (1'h1),
    .RX_PMA_POWER_SAVE (1'b0),
    .RX_PMA_RSV0 (16'h0000),
    .RX_PROGDIV_CFG (0.000000),
    .RX_PROGDIV_RATE (16'h0001),
    .RX_RESLOAD_CTRL (4'b0000),
    .RX_RESLOAD_OVRD (1'b0),
    .RX_SAMPLE_PERIOD (3'b111),
    .RX_SIG_VALID_DLY (11),
    .RX_SUM_DFETAPREP_EN (1'b0),
    .RX_SUM_IREF_TUNE (4'b0100),
    .RX_SUM_RESLOAD_CTRL (4'b0011),
    .RX_SUM_VCMTUNE (4'b0110),
    .RX_SUM_VCM_OVWR (1'b0),
    .RX_SUM_VREF_TUNE (3'b100),
    .RX_TUNE_AFE_OS (2'b00),
    .RX_VREG_CTRL (3'b101),
    .RX_VREG_PDB (1'b1),
    .RX_WIDEMODE_CDR (2'b00),
    .RX_WIDEMODE_CDR_GEN3 (2'b00),
    .RX_WIDEMODE_CDR_GEN4 (2'b01),
    .RX_XCLK_SEL ("RXDES"),
    .RX_XMODE_SEL (1'b0),
    .SAMPLE_CLK_PHASE (1'b0),
    .SAS_12G_MODE (1'b0),
    .SATA_BURST_SEQ_LEN (4'b1111),
    .SATA_BURST_VAL (3'b100),
    .SATA_CPLL_CFG ("VCO_3000MHZ"),
    .SATA_EIDLE_VAL (3'b100),
    .SHOW_REALIGN_COMMA ("TRUE"),
    .SIM_MODE ("FAST"),
    .SIM_RECEIVER_DETECT_PASS ("TRUE"),
    .SIM_RESET_SPEEDUP ("TRUE"),
    .SIM_TX_EIDLE_DRIVE_LEVEL ("Z"),
    .SRSTMODE (1'b0),
    .TAPDLY_SET_TX (2'h0),
    .TEMPERATURE_PAR (4'b0010),
    .TERM_RCAL_CFG (15'b100001000010001),
    .TERM_RCAL_OVRD (3'b000),
    .TRANS_TIME_RATE (8'h0e),
    .TST_RSV0 (8'h00),
    .TST_RSV1 (8'h00),
    .TXBUF_EN ("TRUE"),
    .TXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
    .TXDLY_CFG (16'h8010),
    .TXDLY_LCFG (16'h0030),
    .TXDRVBIAS_N (4'b1010),
    .TXFIFO_ADDR_CFG ("LOW"),
    .TXGBOX_FIFO_INIT_RD_ADDR (4),
    .TXGEARBOX_EN ("FALSE"),
    .TXOUT_DIV (TX_OUT_DIV),
    .TXPCSRESET_TIME (5'b00011),
    .TXPHDLY_CFG0 (16'h6070),
    .TXPHDLY_CFG1 (16'h000f),
    .TXPH_CFG (16'h0323),
    .TXPH_CFG2 (16'h0000),
    .TXPH_MONITOR_SEL (5'b00000),
    .TXPI_CFG (16'h0054),
    .TXPI_CFG0 (2'b00),
    .TXPI_CFG1 (2'b00),
    .TXPI_CFG2 (2'b00),
    .TXPI_CFG3 (1'b0),
    .TXPI_CFG4 (1'b0),
    .TXPI_CFG5 (3'b000),
    .TXPI_GRAY_SEL (1'b0),
    .TXPI_INVSTROBE_SEL (1'b0),
    .TXPI_LPM (1'b0),
    .TXPI_PPM (1'b0),
    .TXPI_PPMCLK_SEL ("TXUSRCLK2"),
    .TXPI_PPM_CFG (8'b00000000),
    .TXPI_SYNFREQ_PPM (3'b001),
    .TXPI_VREFSEL (1'b0),
    .TXPMARESET_TIME (5'b00011),
    .TXREFCLKDIV2_SEL (1'b0),
    .TXSYNC_MULTILANE (1'b1),
    .TXSYNC_OVRD (1'b0),
    .TXSYNC_SKIP_DA (1'b0),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .TX_CLKMUX_EN (1'b1),
    .TX_DATA_WIDTH (40),
    .TX_DCC_LOOP_RST_CFG (16'h0004),
    .TX_DEEMPH0 (6'b000000),
    .TX_DEEMPH1 (6'b000000),
    .TX_DEEMPH2 (6'b000000),
    .TX_DEEMPH3 (6'b000000),
    .TX_DIVRESET_TIME (5'b00001),
    .TX_DRIVE_MODE ("DIRECT"),
    .TX_DRVMUX_CTRL (2),
    .TX_EIDLE_ASSERT_DELAY (3'b100),
    .TX_EIDLE_DEASSERT_DELAY (3'b011),
    .TX_FABINT_USRCLK_FLOP (1'b0),
    .TX_FIFO_BYP_EN (1'b0),
    .TX_IDLE_DATA_ZERO (1'b0),
    .TX_INT_DATAWIDTH (1'h1),
    .TX_LOOPBACK_DRIVE_HIZ ("FALSE"),
    .TX_MAINCURSOR_SEL (1'b0),
    .TX_MARGIN_FULL_0 (7'b1011111),
    .TX_MARGIN_FULL_1 (7'b1011110),
    .TX_MARGIN_FULL_2 (7'b1011100),
    .TX_MARGIN_FULL_3 (7'b1011010),
    .TX_MARGIN_FULL_4 (7'b1011000),
    .TX_MARGIN_LOW_0 (7'b1000110),
    .TX_MARGIN_LOW_1 (7'b1000101),
    .TX_MARGIN_LOW_2 (7'b1000011),
    .TX_MARGIN_LOW_3 (7'b1000010),
    .TX_MARGIN_LOW_4 (7'b1000000),
    .TX_PHICAL_CFG0 (16'h0000),
    .TX_PHICAL_CFG1 (16'h7e00),
    .TX_PHICAL_CFG2 (16'h0201),
    .TX_PI_BIASSET (1'h1),
    .TX_PI_IBIAS_MID (2'b00),
    .TX_PMADATA_OPT (1'b0),
    .TX_PMA_POWER_SAVE (1'b0),
    .TX_PMA_RSV0 (16'h0008),
    .TX_PREDRV_CTRL (2),
    .TX_PROGCLK_SEL ("PREPI"),
    .TX_PROGDIV_CFG (0.000000),
    .TX_PROGDIV_RATE (16'h0001),
    .TX_QPI_STATUS_EN (1'b0),
    .TX_RXDETECT_CFG (14'h0032),
    .TX_RXDETECT_REF (4),
    .TX_SAMPLE_PERIOD (3'b111),
    .TX_SARC_LPBK_ENB (1'b0),
    .TX_SW_MEAS (2'b00),
    .TX_VREG_CTRL (3'b000),
    .TX_VREG_PDB (1'b0),
    .TX_VREG_VREFSEL (2'b00),
    .TX_XCLK_SEL ("TXOUT"),
    .USB_BOTH_BURST_IDLE (1'b0),
    .USB_BURSTMAX_U3WAKE (7'b1111111),
    .USB_BURSTMIN_U3WAKE (7'b1100011),
    .USB_CLK_COR_EQ_EN (1'b0),
    .USB_EXT_CNTL (1'b1),
    .USB_IDLEMAX_POLLING (10'b1010111011),
    .USB_IDLEMIN_POLLING (10'b0100101011),
    .USB_LFPSPING_BURST (9'b000000101),
    .USB_LFPSPOLLING_BURST (9'b000110001),
    .USB_LFPSPOLLING_IDLE_MS (9'b000000100),
    .USB_LFPSU1EXIT_BURST (9'b000011101),
    .USB_LFPSU2LPEXIT_BURST_MS (9'b001100011),
    .USB_LFPSU3WAKE_BURST_MS (9'b111110011),
    .USB_LFPS_TPERIOD (4'b0011),
    .USB_LFPS_TPERIOD_ACCURATE (1'b1),
    .USB_MODE (1'b0),
    .USB_PCIE_ERR_REP_DIS (1'b0),
    .USB_PING_SATA_MAX_INIT (21),
    .USB_PING_SATA_MIN_INIT (12),
    .USB_POLL_SATA_MAX_BURST (8),
    .USB_POLL_SATA_MIN_BURST (4),
    .USB_RAW_ELEC (1'b0),
    .USB_RXIDLE_P0_CTRL (1'b1),
    .USB_TXIDLE_TUNE_ENABLE (1'b1),
    .USB_U1_SATA_MAX_WAKE (7),
    .USB_U1_SATA_MIN_WAKE (4),
    .USB_U2_SAS_MAX_COM (64),
    .USB_U2_SAS_MIN_COM (36),
    .USE_PCS_CLK_PHASE_SEL (1'b0),
    .Y_ALL_MODE (1'b0))
  i_gthe4_channel (
    .BUFGTCE (),
    .BUFGTCEMASK (),
    .BUFGTDIV (),
    .BUFGTRESET (),
    .BUFGTRSTMASK (),
    .CDRSTEPDIR (1'd0),
    .CDRSTEPSQ (1'd0),
    .CDRSTEPSX (1'd0),
    .CFGRESET (1'd0),
    .CLKRSVD0 (1'd0),
    .CLKRSVD1 (1'd0),
    .CPLLFBCLKLOST (),
    .CPLLFREQLOCK (1'd0),
    .CPLLLOCK (cpll_locked_s),
    .CPLLLOCKDETCLK (up_clk),
    .CPLLLOCKEN (1'd1),
    .CPLLPD (1'b0),
    .CPLLREFCLKLOST (),
    .CPLLREFCLKSEL (3'b001),
    .CPLLRESET (up_cpll_rst),
    .DMONFIFORESET (1'd0),
    .DMONITORCLK (1'd0),
    .DMONITOROUT (),
    .DMONITOROUTCLK (),
    .DRPADDR (up_addr_int[9:0]),
    .DRPCLK (up_clk),
    .DRPDI (up_wdata_int),
    .DRPDO (up_rdata_s),
    .DRPEN (up_enb_int),
    .DRPRDY (up_ready_s),
    .DRPRST (1'd0),
    .DRPWE (up_wr_int),
    .EYESCANDATAERROR (),
    .EYESCANRESET (1'd0),
    .EYESCANTRIGGER (1'd0),
    .FREQOS (1'd0),
    .GTGREFCLK (1'd0),
    .GTHRXN (rx_n),
    .GTHRXP (rx_p),
    .GTHTXN (tx_n),
    .GTHTXP (tx_p),
    .GTNORTHREFCLK0 (1'd0),
    .GTNORTHREFCLK1 (1'd0),
    .GTPOWERGOOD (),
    .GTREFCLK0 (cpll_ref_clk),
    .GTREFCLK1 (1'd0),
    .GTREFCLKMONITOR (),
    .GTRSVD (15'd0),
    .GTRXRESET (up_rx_rst),
    .GTRXRESETSEL (1'd0),
    .GTSOUTHREFCLK0 (1'd0),
    .GTSOUTHREFCLK1 (1'd0),
    .GTTXRESET (up_tx_rst),
    .GTTXRESETSEL (1'd0),
    .INCPCTRL (1'd0),
    .LOOPBACK (3'd0),
    .PCIEEQRXEQADAPTDONE (1'd0),
    .PCIERATEGEN3 (),
    .PCIERATEIDLE (),
    .PCIERATEQPLLPD (),
    .PCIERATEQPLLRESET (),
    .PCIERSTIDLE (1'd0),
    .PCIERSTTXSYNCSTART (1'd0),
    .PCIESYNCTXSYNCDONE (),
    .PCIEUSERGEN3RDY (),
    .PCIEUSERPHYSTATUSRST (),
    .PCIEUSERRATEDONE (1'd0),
    .PCIEUSERRATESTART (),
    .PCSRSVDIN (16'd0),
    .PCSRSVDOUT (),
    .PHYSTATUS (),
    .PINRSRVDAS (),
    .POWERPRESENT (),
    .QPLL0CLK (qpll2ch_clk),
    .QPLL0FREQLOCK (1'd0),
    .QPLL0REFCLK (qpll2ch_ref_clk),
    .QPLL1CLK (1'd0),
    .QPLL1FREQLOCK (1'd0),
    .QPLL1REFCLK (1'd0),
    .RESETEXCEPTION (),
    .RESETOVRD (1'd0),
    .RX8B10BEN (1'd1),
    .RXAFECFOKEN (1'b1),
    .RXBUFRESET (1'd0),
    .RXBUFSTATUS (),
    .RXBYTEISALIGNED (),
    .RXBYTEREALIGN (),
    .RXCDRFREQRESET (1'd0),
    .RXCDRHOLD (1'd0),
    .RXCDRLOCK (),
    .RXCDROVRDEN (1'd0),
    .RXCDRPHDONE (),
    .RXCDRRESET (1'd0),
    .RXCHANBONDSEQ (),
    .RXCHANISALIGNED (),
    .RXCHANREALIGN (),
    .RXCHBONDEN (1'd0),
    .RXCHBONDI (5'd0),
    .RXCHBONDLEVEL (3'd0),
    .RXCHBONDMASTER (1'd0),
    .RXCHBONDO (),
    .RXCHBONDSLAVE (1'd0),
    .RXCKCALDONE (),
    .RXCKCALRESET (1'd0),
    .RXCKCALSTART (7'd0),
    .RXCLKCORCNT (),
    .RXCOMINITDET (),
    .RXCOMMADET (),
    .RXCOMMADETEN (1'd1),
    .RXCOMSASDET (),
    .RXCOMWAKEDET (),
    .RXCTRL0 ({rx_charisk_open_s, rx_charisk}),
    .RXCTRL1 ({rx_disperr_open_s, rx_disperr}),
    .RXCTRL2 (),
    .RXCTRL3 ({rx_notintable_open_s, rx_notintable}),
    .RXDATA ({rx_data_open_s, rx_data}),
    .RXDATAEXTENDRSVD (),
    .RXDATAVALID (),
    .RXDFEAGCCTRL (2'b01),
    .RXDFEAGCHOLD (1'd0),
    .RXDFEAGCOVRDEN (1'd0),
    .RXDFECFOKFCNUM (4'b1101),
    .RXDFECFOKFEN (1'd0),
    .RXDFECFOKFPULSE (1'd0),
    .RXDFECFOKHOLD (1'd0),
    .RXDFECFOKOVREN (1'd0),
    .RXDFEKHHOLD (1'd0),
    .RXDFEKHOVRDEN (1'd0),
    .RXDFELFHOLD (1'd0),
    .RXDFELFOVRDEN (1'd0),
    .RXDFELPMRESET (1'd0),
    .RXDFETAP10HOLD (1'd0),
    .RXDFETAP10OVRDEN (1'd0),
    .RXDFETAP11HOLD (1'd0),
    .RXDFETAP11OVRDEN (1'd0),
    .RXDFETAP12HOLD (1'd0),
    .RXDFETAP12OVRDEN (1'd0),
    .RXDFETAP13HOLD (1'd0),
    .RXDFETAP13OVRDEN (1'd0),
    .RXDFETAP14HOLD (1'd0),
    .RXDFETAP14OVRDEN (1'd0),
    .RXDFETAP15HOLD (1'd0),
    .RXDFETAP15OVRDEN (1'd0),
    .RXDFETAP2HOLD (1'd0),
    .RXDFETAP2OVRDEN (1'd0),
    .RXDFETAP3HOLD (1'd0),
    .RXDFETAP3OVRDEN (1'd0),
    .RXDFETAP4HOLD (1'd0),
    .RXDFETAP4OVRDEN (1'd0),
    .RXDFETAP5HOLD (1'd0),
    .RXDFETAP5OVRDEN (1'd0),
    .RXDFETAP6HOLD (1'd0),
    .RXDFETAP6OVRDEN (1'd0),
    .RXDFETAP7HOLD (1'd0),
    .RXDFETAP7OVRDEN (1'd0),
    .RXDFETAP8HOLD (1'd0),
    .RXDFETAP8OVRDEN (1'd0),
    .RXDFETAP9HOLD (1'd0),
    .RXDFETAP9OVRDEN (1'd0),
    .RXDFEUTHOLD (1'd0),
    .RXDFEUTOVRDEN (1'd0),
    .RXDFEVPHOLD (1'd0),
    .RXDFEVPOVRDEN (1'd0),
    .RXDFEXYDEN (1'd1),
    .RXDLYBYPASS (1'd1),
    .RXDLYEN (1'd0),
    .RXDLYOVRDEN (1'd0),
    .RXDLYSRESET (1'd0),
    .RXDLYSRESETDONE (),
    .RXELECIDLE (),
    .RXELECIDLEMODE (2'b11),
    .RXEQTRAINING (1'd0),
    .RXGEARBOXSLIP (1'd0),
    .RXHEADER (),
    .RXHEADERVALID (),
    .RXLATCLK (1'd0),
    .RXLFPSTRESETDET (),
    .RXLFPSU2LPEXITDET (),
    .RXLFPSU3WAKEDET (),
    .RXLPMEN (up_rx_lpm_dfe_n),
    .RXLPMGCHOLD (1'd0),
    .RXLPMGCOVRDEN (1'd0),
    .RXLPMHFHOLD (1'd0),
    .RXLPMHFOVRDEN (1'd0),
    .RXLPMLFHOLD (1'd0),
    .RXLPMLFKLOVRDEN (1'd0),
    .RXLPMOSHOLD (1'd0),
    .RXLPMOSOVRDEN (1'd0),
    .RXMCOMMAALIGNEN (rx_calign),
    .RXMONITOROUT (),
    .RXMONITORSEL (2'd0),
    .RXOOBRESET (1'd0),
    .RXOSCALRESET (1'd0),
    .RXOSHOLD (1'd0),
    .RXOSINTDONE (),
    .RXOSINTSTARTED (),
    .RXOSINTSTROBEDONE (),
    .RXOSINTSTROBESTARTED (),
    .RXOSOVRDEN (1'd0),
    .RXOUTCLK (rx_out_clk_s),
    .RXOUTCLKFABRIC (),
    .RXOUTCLKPCS (),
    .RXOUTCLKSEL (up_rx_out_clk_sel),
    .RXPCOMMAALIGNEN (rx_calign),
    .RXPCSRESET (1'd0),
    .RXPD (2'd0),
    .RXPHALIGN (1'd0),
    .RXPHALIGNDONE (),
    .RXPHALIGNEN (1'd0),
    .RXPHALIGNERR (),
    .RXPHDLYPD (1'd1),
    .RXPHDLYRESET (1'd0),
    .RXPHOVRDEN (1'd0),
    .RXPLLCLKSEL (rx_pll_clk_sel_s),
    .RXPMARESET (1'd0),
    .RXPMARESETDONE (),
    .RXPOLARITY (1'd0),
    .RXPRBSCNTRESET (1'd0),
    .RXPRBSERR (),
    .RXPRBSLOCKED (),
    .RXPRBSSEL (4'd0),
    .RXPRGDIVRESETDONE (),
    .RXPROGDIVRESET (1'd0),
    .RXQPIEN (1'd0),
    .RXQPISENN (),
    .RXQPISENP (),
    .RXRATE (rx_rate_m2),
    .RXRATEDONE (),
    .RXRATEMODE (1'd0),
    .RXRECCLKOUT (),
    .RXRESETDONE (rx_rst_done_s),
    .RXSLIDE (1'd0),
    .RXSLIDERDY (),
    .RXSLIPDONE (),
    .RXSLIPOUTCLK (1'd0),
    .RXSLIPOUTCLKRDY (),
    .RXSLIPPMA (1'd0),
    .RXSLIPPMARDY (),
    .RXSTARTOFSEQ (),
    .RXSTATUS (),
    .RXSYNCALLIN (1'd0),
    .RXSYNCDONE (),
    .RXSYNCIN (1'd0),
    .RXSYNCMODE (1'd0),
    .RXSYNCOUT (),
    .RXSYSCLKSEL (rx_sys_clk_sel_s),
    .RXTERMINATION (1'd0),
    .RXUSERRDY (up_rx_user_ready),
    .RXUSRCLK (rx_clk),
    .RXUSRCLK2 (rx_clk),
    .RXVALID (),
    .SIGVALIDCLK (1'd0),
    .TSTIN (20'd0),
    .TX8B10BBYPASS (8'd0),
    .TX8B10BEN (1'd1),
    .TXBUFSTATUS (),
    .TXCOMFINISH (),
    .TXCOMINIT (1'd0),
    .TXCOMSAS (1'd0),
    .TXCOMWAKE (1'd0),
    .TXCTRL0 (16'd0),
    .TXCTRL1 (16'd0),
    .TXCTRL2 ({4'd0, tx_charisk}),
    .TXDATA ({96'd0, tx_data}),
    .TXDATAEXTENDRSVD (8'd0),
    .TXDCCDONE (),
    .TXDCCFORCESTART (1'd0),
    .TXDCCRESET (1'd0),
    .TXDEEMPH (2'd0),
    .TXDETECTRX (1'd0),
    .TXDIFFCTRL (5'b00000),
    .TXDLYBYPASS (1'd1),
    .TXDLYEN (1'd0),
    .TXDLYHOLD (1'd0),
    .TXDLYOVRDEN (1'd0),
    .TXDLYSRESET (1'd0),
    .TXDLYSRESETDONE (),
    .TXDLYUPDOWN (1'd0),
    .TXELECIDLE (1'd0),
    .TXHEADER (6'd0),
    .TXINHIBIT (1'd0),
    .TXLATCLK (1'd0),
    .TXLFPSTRESET (1'd0),
    .TXLFPSU2LPEXIT (1'd0),
    .TXLFPSU3WAKE (1'd0),
    .TXMAINCURSOR (7'b1000000),
    .TXMARGIN (3'd0),
    .TXMUXDCDEXHOLD (1'd0),
    .TXMUXDCDORWREN (1'd0),
    .TXONESZEROS (1'd0),
    .TXOUTCLK (tx_out_clk_s),
    .TXOUTCLKFABRIC (),
    .TXOUTCLKPCS (),
    .TXOUTCLKSEL (up_tx_out_clk_sel),
    .TXPCSRESET (1'd0),
    .TXPD (2'd0),
    .TXPDELECIDLEMODE (1'd0),
    .TXPHALIGN (1'd0),
    .TXPHALIGNDONE (),
    .TXPHALIGNEN (1'd0),
    .TXPHDLYPD (1'd1),
    .TXPHDLYRESET (1'd0),
    .TXPHDLYTSTCLK (1'd0),
    .TXPHINIT (1'd0),
    .TXPHINITDONE (),
    .TXPHOVRDEN (1'd0),
    .TXPIPPMEN (1'd0),
    .TXPIPPMOVRDEN (1'd0),
    .TXPIPPMPD (1'd0),
    .TXPIPPMSEL (1'd0),
    .TXPIPPMSTEPSIZE (5'd0),
    .TXPISOPD (1'd0),
    .TXPLLCLKSEL (tx_pll_clk_sel_s),
    .TXPMARESET (1'd0),
    .TXPMARESETDONE (),
    .TXPOLARITY (1'd0),
    .TXPOSTCURSOR (5'd0),
    .TXPRBSFORCEERR (1'd0),
    .TXPRBSSEL (4'd0),
    .TXPRECURSOR (5'd0),
    .TXPRGDIVRESETDONE (),
    .TXPROGDIVRESET (up_tx_rst),
    .TXQPIBIASEN (1'd0),
    .TXQPISENN (),
    .TXQPISENP (),
    .TXQPIWEAKPUP (1'd0),
    .TXRATE (tx_rate_m2),
    .TXRATEDONE (),
    .TXRATEMODE (1'd0),
    .TXRESETDONE (tx_rst_done_s),
    .TXSEQUENCE (7'd0),
    .TXSWING (1'd0),
    .TXSYNCALLIN (1'd0),
    .TXSYNCDONE (),
    .TXSYNCIN (1'd0),
    .TXSYNCMODE (1'd0),
    .TXSYNCOUT (),
    .TXSYSCLKSEL (tx_sys_clk_sel_s),
    .TXUSERRDY (up_tx_user_ready),
    .TXUSRCLK (tx_clk),
    .TXUSRCLK2 (tx_clk));
  end
  endgenerate

endmodule

// ***************************************************************************
// ***************************************************************************


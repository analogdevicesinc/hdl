// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************
// AUTO GENERATED BY util_adxcvr.pl, DO NOT MODIFY!

`timescale 1ns/1ps

module util_adxcvr #(

  // gtxe2(0), gthe3(1), gthe4(2)

  parameter   integer XCVR_TYPE = 0,

  // qpll-configuration

  parameter   integer QPLL_REFCLK_DIV = 1,
  parameter   integer QPLL_FBDIV_RATIO = 1,
  parameter   [26:0]  QPLL_CFG = 27'h0680181,
  parameter   [ 9:0]  QPLL_FBDIV =  10'b0000110000,

  // cpll-configuration

  parameter   integer CPLL_FBDIV = 2,
  parameter   integer CPLL_FBDIV_4_5 = 5,

  // tx-configuration

  parameter   integer TX_NUM_OF_LANES = 8,
  parameter   integer TX_OUT_DIV = 1,
  parameter   integer TX_CLK25_DIV = 20,

  // rx-configuration

  parameter   integer RX_NUM_OF_LANES = 8,
  parameter   integer RX_OUT_DIV = 1,
  parameter   integer RX_CLK25_DIV = 20,
  parameter   [15:0]  RX_DFE_LPM_CFG = 16'h0104,
  parameter   [31:0]  RX_PMA_CFG = 32'h001e7080,
  parameter   [72:0]  RX_CDR_CFG = 72'h0b000023ff10400020) (

  input           up_rstn,
  input           up_clk,

  input           qpll_ref_clk_0,
  input           up_qpll_rst_0,
  input           cpll_ref_clk_0,
  input           up_cpll_rst_0,

  input           rx_0_p,
  input           rx_0_n,
  output          rx_out_clk_0,
  input           rx_clk_0,
  output  [ 3:0]  rx_charisk_0,
  output  [ 3:0]  rx_disperr_0,
  output  [ 3:0]  rx_notintable_0,
  output  [31:0]  rx_data_0,
  input           rx_calign_0,

  output          tx_0_p,
  output          tx_0_n,
  output          tx_out_clk_0,
  input           tx_clk_0,
  input   [ 3:0]  tx_charisk_0,
  input   [31:0]  tx_data_0,

  input   [ 7:0]  up_cm_sel_0,
  input           up_cm_enb_0,
  input   [11:0]  up_cm_addr_0,
  input           up_cm_wr_0,
  input   [15:0]  up_cm_wdata_0,
  output  [15:0]  up_cm_rdata_0,
  output          up_cm_ready_0,
  input   [ 7:0]  up_es_sel_0,
  input           up_es_enb_0,
  input   [11:0]  up_es_addr_0,
  input           up_es_wr_0,
  input   [15:0]  up_es_wdata_0,
  output  [15:0]  up_es_rdata_0,
  output          up_es_ready_0,
  output          up_rx_pll_locked_0,
  input           up_rx_rst_0,
  input           up_rx_user_ready_0,
  output          up_rx_rst_done_0,
  input           up_rx_lpm_dfe_n_0,
  input   [ 2:0]  up_rx_rate_0,
  input   [ 1:0]  up_rx_sys_clk_sel_0,
  input   [ 2:0]  up_rx_out_clk_sel_0,
  input   [ 7:0]  up_rx_sel_0,
  input           up_rx_enb_0,
  input   [11:0]  up_rx_addr_0,
  input           up_rx_wr_0,
  input   [15:0]  up_rx_wdata_0,
  output  [15:0]  up_rx_rdata_0,
  output          up_rx_ready_0,
  output          up_tx_pll_locked_0,
  input           up_tx_rst_0,
  input           up_tx_user_ready_0,
  output          up_tx_rst_done_0,
  input           up_tx_lpm_dfe_n_0,
  input   [ 2:0]  up_tx_rate_0,
  input   [ 1:0]  up_tx_sys_clk_sel_0,
  input   [ 2:0]  up_tx_out_clk_sel_0,
  input   [ 7:0]  up_tx_sel_0,
  input           up_tx_enb_0,
  input   [11:0]  up_tx_addr_0,
  input           up_tx_wr_0,
  input   [15:0]  up_tx_wdata_0,
  output  [15:0]  up_tx_rdata_0,
  output          up_tx_ready_0,

  input           cpll_ref_clk_1,
  input           up_cpll_rst_1,

  input           rx_1_p,
  input           rx_1_n,
  output          rx_out_clk_1,
  input           rx_clk_1,
  output  [ 3:0]  rx_charisk_1,
  output  [ 3:0]  rx_disperr_1,
  output  [ 3:0]  rx_notintable_1,
  output  [31:0]  rx_data_1,
  input           rx_calign_1,

  output          tx_1_p,
  output          tx_1_n,
  output          tx_out_clk_1,
  input           tx_clk_1,
  input   [ 3:0]  tx_charisk_1,
  input   [31:0]  tx_data_1,

  input   [ 7:0]  up_es_sel_1,
  input           up_es_enb_1,
  input   [11:0]  up_es_addr_1,
  input           up_es_wr_1,
  input   [15:0]  up_es_wdata_1,
  output  [15:0]  up_es_rdata_1,
  output          up_es_ready_1,
  output          up_rx_pll_locked_1,
  input           up_rx_rst_1,
  input           up_rx_user_ready_1,
  output          up_rx_rst_done_1,
  input           up_rx_lpm_dfe_n_1,
  input   [ 2:0]  up_rx_rate_1,
  input   [ 1:0]  up_rx_sys_clk_sel_1,
  input   [ 2:0]  up_rx_out_clk_sel_1,
  input   [ 7:0]  up_rx_sel_1,
  input           up_rx_enb_1,
  input   [11:0]  up_rx_addr_1,
  input           up_rx_wr_1,
  input   [15:0]  up_rx_wdata_1,
  output  [15:0]  up_rx_rdata_1,
  output          up_rx_ready_1,
  output          up_tx_pll_locked_1,
  input           up_tx_rst_1,
  input           up_tx_user_ready_1,
  output          up_tx_rst_done_1,
  input           up_tx_lpm_dfe_n_1,
  input   [ 2:0]  up_tx_rate_1,
  input   [ 1:0]  up_tx_sys_clk_sel_1,
  input   [ 2:0]  up_tx_out_clk_sel_1,
  input   [ 7:0]  up_tx_sel_1,
  input           up_tx_enb_1,
  input   [11:0]  up_tx_addr_1,
  input           up_tx_wr_1,
  input   [15:0]  up_tx_wdata_1,
  output  [15:0]  up_tx_rdata_1,
  output          up_tx_ready_1,

  input           cpll_ref_clk_2,
  input           up_cpll_rst_2,

  input           rx_2_p,
  input           rx_2_n,
  output          rx_out_clk_2,
  input           rx_clk_2,
  output  [ 3:0]  rx_charisk_2,
  output  [ 3:0]  rx_disperr_2,
  output  [ 3:0]  rx_notintable_2,
  output  [31:0]  rx_data_2,
  input           rx_calign_2,

  output          tx_2_p,
  output          tx_2_n,
  output          tx_out_clk_2,
  input           tx_clk_2,
  input   [ 3:0]  tx_charisk_2,
  input   [31:0]  tx_data_2,

  input   [ 7:0]  up_es_sel_2,
  input           up_es_enb_2,
  input   [11:0]  up_es_addr_2,
  input           up_es_wr_2,
  input   [15:0]  up_es_wdata_2,
  output  [15:0]  up_es_rdata_2,
  output          up_es_ready_2,
  output          up_rx_pll_locked_2,
  input           up_rx_rst_2,
  input           up_rx_user_ready_2,
  output          up_rx_rst_done_2,
  input           up_rx_lpm_dfe_n_2,
  input   [ 2:0]  up_rx_rate_2,
  input   [ 1:0]  up_rx_sys_clk_sel_2,
  input   [ 2:0]  up_rx_out_clk_sel_2,
  input   [ 7:0]  up_rx_sel_2,
  input           up_rx_enb_2,
  input   [11:0]  up_rx_addr_2,
  input           up_rx_wr_2,
  input   [15:0]  up_rx_wdata_2,
  output  [15:0]  up_rx_rdata_2,
  output          up_rx_ready_2,
  output          up_tx_pll_locked_2,
  input           up_tx_rst_2,
  input           up_tx_user_ready_2,
  output          up_tx_rst_done_2,
  input           up_tx_lpm_dfe_n_2,
  input   [ 2:0]  up_tx_rate_2,
  input   [ 1:0]  up_tx_sys_clk_sel_2,
  input   [ 2:0]  up_tx_out_clk_sel_2,
  input   [ 7:0]  up_tx_sel_2,
  input           up_tx_enb_2,
  input   [11:0]  up_tx_addr_2,
  input           up_tx_wr_2,
  input   [15:0]  up_tx_wdata_2,
  output  [15:0]  up_tx_rdata_2,
  output          up_tx_ready_2,

  input           cpll_ref_clk_3,
  input           up_cpll_rst_3,

  input           rx_3_p,
  input           rx_3_n,
  output          rx_out_clk_3,
  input           rx_clk_3,
  output  [ 3:0]  rx_charisk_3,
  output  [ 3:0]  rx_disperr_3,
  output  [ 3:0]  rx_notintable_3,
  output  [31:0]  rx_data_3,
  input           rx_calign_3,

  output          tx_3_p,
  output          tx_3_n,
  output          tx_out_clk_3,
  input           tx_clk_3,
  input   [ 3:0]  tx_charisk_3,
  input   [31:0]  tx_data_3,

  input   [ 7:0]  up_es_sel_3,
  input           up_es_enb_3,
  input   [11:0]  up_es_addr_3,
  input           up_es_wr_3,
  input   [15:0]  up_es_wdata_3,
  output  [15:0]  up_es_rdata_3,
  output          up_es_ready_3,
  output          up_rx_pll_locked_3,
  input           up_rx_rst_3,
  input           up_rx_user_ready_3,
  output          up_rx_rst_done_3,
  input           up_rx_lpm_dfe_n_3,
  input   [ 2:0]  up_rx_rate_3,
  input   [ 1:0]  up_rx_sys_clk_sel_3,
  input   [ 2:0]  up_rx_out_clk_sel_3,
  input   [ 7:0]  up_rx_sel_3,
  input           up_rx_enb_3,
  input   [11:0]  up_rx_addr_3,
  input           up_rx_wr_3,
  input   [15:0]  up_rx_wdata_3,
  output  [15:0]  up_rx_rdata_3,
  output          up_rx_ready_3,
  output          up_tx_pll_locked_3,
  input           up_tx_rst_3,
  input           up_tx_user_ready_3,
  output          up_tx_rst_done_3,
  input           up_tx_lpm_dfe_n_3,
  input   [ 2:0]  up_tx_rate_3,
  input   [ 1:0]  up_tx_sys_clk_sel_3,
  input   [ 2:0]  up_tx_out_clk_sel_3,
  input   [ 7:0]  up_tx_sel_3,
  input           up_tx_enb_3,
  input   [11:0]  up_tx_addr_3,
  input           up_tx_wr_3,
  input   [15:0]  up_tx_wdata_3,
  output  [15:0]  up_tx_rdata_3,
  output          up_tx_ready_3,

  input           qpll_ref_clk_4,
  input           up_qpll_rst_4,
  input           cpll_ref_clk_4,
  input           up_cpll_rst_4,

  input           rx_4_p,
  input           rx_4_n,
  output          rx_out_clk_4,
  input           rx_clk_4,
  output  [ 3:0]  rx_charisk_4,
  output  [ 3:0]  rx_disperr_4,
  output  [ 3:0]  rx_notintable_4,
  output  [31:0]  rx_data_4,
  input           rx_calign_4,

  output          tx_4_p,
  output          tx_4_n,
  output          tx_out_clk_4,
  input           tx_clk_4,
  input   [ 3:0]  tx_charisk_4,
  input   [31:0]  tx_data_4,

  input   [ 7:0]  up_cm_sel_4,
  input           up_cm_enb_4,
  input   [11:0]  up_cm_addr_4,
  input           up_cm_wr_4,
  input   [15:0]  up_cm_wdata_4,
  output  [15:0]  up_cm_rdata_4,
  output          up_cm_ready_4,
  input   [ 7:0]  up_es_sel_4,
  input           up_es_enb_4,
  input   [11:0]  up_es_addr_4,
  input           up_es_wr_4,
  input   [15:0]  up_es_wdata_4,
  output  [15:0]  up_es_rdata_4,
  output          up_es_ready_4,
  output          up_rx_pll_locked_4,
  input           up_rx_rst_4,
  input           up_rx_user_ready_4,
  output          up_rx_rst_done_4,
  input           up_rx_lpm_dfe_n_4,
  input   [ 2:0]  up_rx_rate_4,
  input   [ 1:0]  up_rx_sys_clk_sel_4,
  input   [ 2:0]  up_rx_out_clk_sel_4,
  input   [ 7:0]  up_rx_sel_4,
  input           up_rx_enb_4,
  input   [11:0]  up_rx_addr_4,
  input           up_rx_wr_4,
  input   [15:0]  up_rx_wdata_4,
  output  [15:0]  up_rx_rdata_4,
  output          up_rx_ready_4,
  output          up_tx_pll_locked_4,
  input           up_tx_rst_4,
  input           up_tx_user_ready_4,
  output          up_tx_rst_done_4,
  input           up_tx_lpm_dfe_n_4,
  input   [ 2:0]  up_tx_rate_4,
  input   [ 1:0]  up_tx_sys_clk_sel_4,
  input   [ 2:0]  up_tx_out_clk_sel_4,
  input   [ 7:0]  up_tx_sel_4,
  input           up_tx_enb_4,
  input   [11:0]  up_tx_addr_4,
  input           up_tx_wr_4,
  input   [15:0]  up_tx_wdata_4,
  output  [15:0]  up_tx_rdata_4,
  output          up_tx_ready_4,

  input           cpll_ref_clk_5,
  input           up_cpll_rst_5,

  input           rx_5_p,
  input           rx_5_n,
  output          rx_out_clk_5,
  input           rx_clk_5,
  output  [ 3:0]  rx_charisk_5,
  output  [ 3:0]  rx_disperr_5,
  output  [ 3:0]  rx_notintable_5,
  output  [31:0]  rx_data_5,
  input           rx_calign_5,

  output          tx_5_p,
  output          tx_5_n,
  output          tx_out_clk_5,
  input           tx_clk_5,
  input   [ 3:0]  tx_charisk_5,
  input   [31:0]  tx_data_5,

  input   [ 7:0]  up_es_sel_5,
  input           up_es_enb_5,
  input   [11:0]  up_es_addr_5,
  input           up_es_wr_5,
  input   [15:0]  up_es_wdata_5,
  output  [15:0]  up_es_rdata_5,
  output          up_es_ready_5,
  output          up_rx_pll_locked_5,
  input           up_rx_rst_5,
  input           up_rx_user_ready_5,
  output          up_rx_rst_done_5,
  input           up_rx_lpm_dfe_n_5,
  input   [ 2:0]  up_rx_rate_5,
  input   [ 1:0]  up_rx_sys_clk_sel_5,
  input   [ 2:0]  up_rx_out_clk_sel_5,
  input   [ 7:0]  up_rx_sel_5,
  input           up_rx_enb_5,
  input   [11:0]  up_rx_addr_5,
  input           up_rx_wr_5,
  input   [15:0]  up_rx_wdata_5,
  output  [15:0]  up_rx_rdata_5,
  output          up_rx_ready_5,
  output          up_tx_pll_locked_5,
  input           up_tx_rst_5,
  input           up_tx_user_ready_5,
  output          up_tx_rst_done_5,
  input           up_tx_lpm_dfe_n_5,
  input   [ 2:0]  up_tx_rate_5,
  input   [ 1:0]  up_tx_sys_clk_sel_5,
  input   [ 2:0]  up_tx_out_clk_sel_5,
  input   [ 7:0]  up_tx_sel_5,
  input           up_tx_enb_5,
  input   [11:0]  up_tx_addr_5,
  input           up_tx_wr_5,
  input   [15:0]  up_tx_wdata_5,
  output  [15:0]  up_tx_rdata_5,
  output          up_tx_ready_5,

  input           cpll_ref_clk_6,
  input           up_cpll_rst_6,

  input           rx_6_p,
  input           rx_6_n,
  output          rx_out_clk_6,
  input           rx_clk_6,
  output  [ 3:0]  rx_charisk_6,
  output  [ 3:0]  rx_disperr_6,
  output  [ 3:0]  rx_notintable_6,
  output  [31:0]  rx_data_6,
  input           rx_calign_6,

  output          tx_6_p,
  output          tx_6_n,
  output          tx_out_clk_6,
  input           tx_clk_6,
  input   [ 3:0]  tx_charisk_6,
  input   [31:0]  tx_data_6,

  input   [ 7:0]  up_es_sel_6,
  input           up_es_enb_6,
  input   [11:0]  up_es_addr_6,
  input           up_es_wr_6,
  input   [15:0]  up_es_wdata_6,
  output  [15:0]  up_es_rdata_6,
  output          up_es_ready_6,
  output          up_rx_pll_locked_6,
  input           up_rx_rst_6,
  input           up_rx_user_ready_6,
  output          up_rx_rst_done_6,
  input           up_rx_lpm_dfe_n_6,
  input   [ 2:0]  up_rx_rate_6,
  input   [ 1:0]  up_rx_sys_clk_sel_6,
  input   [ 2:0]  up_rx_out_clk_sel_6,
  input   [ 7:0]  up_rx_sel_6,
  input           up_rx_enb_6,
  input   [11:0]  up_rx_addr_6,
  input           up_rx_wr_6,
  input   [15:0]  up_rx_wdata_6,
  output  [15:0]  up_rx_rdata_6,
  output          up_rx_ready_6,
  output          up_tx_pll_locked_6,
  input           up_tx_rst_6,
  input           up_tx_user_ready_6,
  output          up_tx_rst_done_6,
  input           up_tx_lpm_dfe_n_6,
  input   [ 2:0]  up_tx_rate_6,
  input   [ 1:0]  up_tx_sys_clk_sel_6,
  input   [ 2:0]  up_tx_out_clk_sel_6,
  input   [ 7:0]  up_tx_sel_6,
  input           up_tx_enb_6,
  input   [11:0]  up_tx_addr_6,
  input           up_tx_wr_6,
  input   [15:0]  up_tx_wdata_6,
  output  [15:0]  up_tx_rdata_6,
  output          up_tx_ready_6,

  input           cpll_ref_clk_7,
  input           up_cpll_rst_7,

  input           rx_7_p,
  input           rx_7_n,
  output          rx_out_clk_7,
  input           rx_clk_7,
  output  [ 3:0]  rx_charisk_7,
  output  [ 3:0]  rx_disperr_7,
  output  [ 3:0]  rx_notintable_7,
  output  [31:0]  rx_data_7,
  input           rx_calign_7,

  output          tx_7_p,
  output          tx_7_n,
  output          tx_out_clk_7,
  input           tx_clk_7,
  input   [ 3:0]  tx_charisk_7,
  input   [31:0]  tx_data_7,

  input   [ 7:0]  up_es_sel_7,
  input           up_es_enb_7,
  input   [11:0]  up_es_addr_7,
  input           up_es_wr_7,
  input   [15:0]  up_es_wdata_7,
  output  [15:0]  up_es_rdata_7,
  output          up_es_ready_7,
  output          up_rx_pll_locked_7,
  input           up_rx_rst_7,
  input           up_rx_user_ready_7,
  output          up_rx_rst_done_7,
  input           up_rx_lpm_dfe_n_7,
  input   [ 2:0]  up_rx_rate_7,
  input   [ 1:0]  up_rx_sys_clk_sel_7,
  input   [ 2:0]  up_rx_out_clk_sel_7,
  input   [ 7:0]  up_rx_sel_7,
  input           up_rx_enb_7,
  input   [11:0]  up_rx_addr_7,
  input           up_rx_wr_7,
  input   [15:0]  up_rx_wdata_7,
  output  [15:0]  up_rx_rdata_7,
  output          up_rx_ready_7,
  output          up_tx_pll_locked_7,
  input           up_tx_rst_7,
  input           up_tx_user_ready_7,
  output          up_tx_rst_done_7,
  input           up_tx_lpm_dfe_n_7,
  input   [ 2:0]  up_tx_rate_7,
  input   [ 1:0]  up_tx_sys_clk_sel_7,
  input   [ 2:0]  up_tx_out_clk_sel_7,
  input   [ 7:0]  up_tx_sel_7,
  input           up_tx_enb_7,
  input   [11:0]  up_tx_addr_7,
  input           up_tx_wr_7,
  input   [15:0]  up_tx_wdata_7,
  output  [15:0]  up_tx_rdata_7,
  output          up_tx_ready_7,

  input           qpll_ref_clk_8,
  input           up_qpll_rst_8,
  input           cpll_ref_clk_8,
  input           up_cpll_rst_8,

  input           rx_8_p,
  input           rx_8_n,
  output          rx_out_clk_8,
  input           rx_clk_8,
  output  [ 3:0]  rx_charisk_8,
  output  [ 3:0]  rx_disperr_8,
  output  [ 3:0]  rx_notintable_8,
  output  [31:0]  rx_data_8,
  input           rx_calign_8,

  output          tx_8_p,
  output          tx_8_n,
  output          tx_out_clk_8,
  input           tx_clk_8,
  input   [ 3:0]  tx_charisk_8,
  input   [31:0]  tx_data_8,

  input   [ 7:0]  up_cm_sel_8,
  input           up_cm_enb_8,
  input   [11:0]  up_cm_addr_8,
  input           up_cm_wr_8,
  input   [15:0]  up_cm_wdata_8,
  output  [15:0]  up_cm_rdata_8,
  output          up_cm_ready_8,
  input   [ 7:0]  up_es_sel_8,
  input           up_es_enb_8,
  input   [11:0]  up_es_addr_8,
  input           up_es_wr_8,
  input   [15:0]  up_es_wdata_8,
  output  [15:0]  up_es_rdata_8,
  output          up_es_ready_8,
  output          up_rx_pll_locked_8,
  input           up_rx_rst_8,
  input           up_rx_user_ready_8,
  output          up_rx_rst_done_8,
  input           up_rx_lpm_dfe_n_8,
  input   [ 2:0]  up_rx_rate_8,
  input   [ 1:0]  up_rx_sys_clk_sel_8,
  input   [ 2:0]  up_rx_out_clk_sel_8,
  input   [ 7:0]  up_rx_sel_8,
  input           up_rx_enb_8,
  input   [11:0]  up_rx_addr_8,
  input           up_rx_wr_8,
  input   [15:0]  up_rx_wdata_8,
  output  [15:0]  up_rx_rdata_8,
  output          up_rx_ready_8,
  output          up_tx_pll_locked_8,
  input           up_tx_rst_8,
  input           up_tx_user_ready_8,
  output          up_tx_rst_done_8,
  input           up_tx_lpm_dfe_n_8,
  input   [ 2:0]  up_tx_rate_8,
  input   [ 1:0]  up_tx_sys_clk_sel_8,
  input   [ 2:0]  up_tx_out_clk_sel_8,
  input   [ 7:0]  up_tx_sel_8,
  input           up_tx_enb_8,
  input   [11:0]  up_tx_addr_8,
  input           up_tx_wr_8,
  input   [15:0]  up_tx_wdata_8,
  output  [15:0]  up_tx_rdata_8,
  output          up_tx_ready_8,

  input           cpll_ref_clk_9,
  input           up_cpll_rst_9,

  input           rx_9_p,
  input           rx_9_n,
  output          rx_out_clk_9,
  input           rx_clk_9,
  output  [ 3:0]  rx_charisk_9,
  output  [ 3:0]  rx_disperr_9,
  output  [ 3:0]  rx_notintable_9,
  output  [31:0]  rx_data_9,
  input           rx_calign_9,

  output          tx_9_p,
  output          tx_9_n,
  output          tx_out_clk_9,
  input           tx_clk_9,
  input   [ 3:0]  tx_charisk_9,
  input   [31:0]  tx_data_9,

  input   [ 7:0]  up_es_sel_9,
  input           up_es_enb_9,
  input   [11:0]  up_es_addr_9,
  input           up_es_wr_9,
  input   [15:0]  up_es_wdata_9,
  output  [15:0]  up_es_rdata_9,
  output          up_es_ready_9,
  output          up_rx_pll_locked_9,
  input           up_rx_rst_9,
  input           up_rx_user_ready_9,
  output          up_rx_rst_done_9,
  input           up_rx_lpm_dfe_n_9,
  input   [ 2:0]  up_rx_rate_9,
  input   [ 1:0]  up_rx_sys_clk_sel_9,
  input   [ 2:0]  up_rx_out_clk_sel_9,
  input   [ 7:0]  up_rx_sel_9,
  input           up_rx_enb_9,
  input   [11:0]  up_rx_addr_9,
  input           up_rx_wr_9,
  input   [15:0]  up_rx_wdata_9,
  output  [15:0]  up_rx_rdata_9,
  output          up_rx_ready_9,
  output          up_tx_pll_locked_9,
  input           up_tx_rst_9,
  input           up_tx_user_ready_9,
  output          up_tx_rst_done_9,
  input           up_tx_lpm_dfe_n_9,
  input   [ 2:0]  up_tx_rate_9,
  input   [ 1:0]  up_tx_sys_clk_sel_9,
  input   [ 2:0]  up_tx_out_clk_sel_9,
  input   [ 7:0]  up_tx_sel_9,
  input           up_tx_enb_9,
  input   [11:0]  up_tx_addr_9,
  input           up_tx_wr_9,
  input   [15:0]  up_tx_wdata_9,
  output  [15:0]  up_tx_rdata_9,
  output          up_tx_ready_9,

  input           cpll_ref_clk_10,
  input           up_cpll_rst_10,

  input           rx_10_p,
  input           rx_10_n,
  output          rx_out_clk_10,
  input           rx_clk_10,
  output  [ 3:0]  rx_charisk_10,
  output  [ 3:0]  rx_disperr_10,
  output  [ 3:0]  rx_notintable_10,
  output  [31:0]  rx_data_10,
  input           rx_calign_10,

  output          tx_10_p,
  output          tx_10_n,
  output          tx_out_clk_10,
  input           tx_clk_10,
  input   [ 3:0]  tx_charisk_10,
  input   [31:0]  tx_data_10,

  input   [ 7:0]  up_es_sel_10,
  input           up_es_enb_10,
  input   [11:0]  up_es_addr_10,
  input           up_es_wr_10,
  input   [15:0]  up_es_wdata_10,
  output  [15:0]  up_es_rdata_10,
  output          up_es_ready_10,
  output          up_rx_pll_locked_10,
  input           up_rx_rst_10,
  input           up_rx_user_ready_10,
  output          up_rx_rst_done_10,
  input           up_rx_lpm_dfe_n_10,
  input   [ 2:0]  up_rx_rate_10,
  input   [ 1:0]  up_rx_sys_clk_sel_10,
  input   [ 2:0]  up_rx_out_clk_sel_10,
  input   [ 7:0]  up_rx_sel_10,
  input           up_rx_enb_10,
  input   [11:0]  up_rx_addr_10,
  input           up_rx_wr_10,
  input   [15:0]  up_rx_wdata_10,
  output  [15:0]  up_rx_rdata_10,
  output          up_rx_ready_10,
  output          up_tx_pll_locked_10,
  input           up_tx_rst_10,
  input           up_tx_user_ready_10,
  output          up_tx_rst_done_10,
  input           up_tx_lpm_dfe_n_10,
  input   [ 2:0]  up_tx_rate_10,
  input   [ 1:0]  up_tx_sys_clk_sel_10,
  input   [ 2:0]  up_tx_out_clk_sel_10,
  input   [ 7:0]  up_tx_sel_10,
  input           up_tx_enb_10,
  input   [11:0]  up_tx_addr_10,
  input           up_tx_wr_10,
  input   [15:0]  up_tx_wdata_10,
  output  [15:0]  up_tx_rdata_10,
  output          up_tx_ready_10,

  input           cpll_ref_clk_11,
  input           up_cpll_rst_11,

  input           rx_11_p,
  input           rx_11_n,
  output          rx_out_clk_11,
  input           rx_clk_11,
  output  [ 3:0]  rx_charisk_11,
  output  [ 3:0]  rx_disperr_11,
  output  [ 3:0]  rx_notintable_11,
  output  [31:0]  rx_data_11,
  input           rx_calign_11,

  output          tx_11_p,
  output          tx_11_n,
  output          tx_out_clk_11,
  input           tx_clk_11,
  input   [ 3:0]  tx_charisk_11,
  input   [31:0]  tx_data_11,

  input   [ 7:0]  up_es_sel_11,
  input           up_es_enb_11,
  input   [11:0]  up_es_addr_11,
  input           up_es_wr_11,
  input   [15:0]  up_es_wdata_11,
  output  [15:0]  up_es_rdata_11,
  output          up_es_ready_11,
  output          up_rx_pll_locked_11,
  input           up_rx_rst_11,
  input           up_rx_user_ready_11,
  output          up_rx_rst_done_11,
  input           up_rx_lpm_dfe_n_11,
  input   [ 2:0]  up_rx_rate_11,
  input   [ 1:0]  up_rx_sys_clk_sel_11,
  input   [ 2:0]  up_rx_out_clk_sel_11,
  input   [ 7:0]  up_rx_sel_11,
  input           up_rx_enb_11,
  input   [11:0]  up_rx_addr_11,
  input           up_rx_wr_11,
  input   [15:0]  up_rx_wdata_11,
  output  [15:0]  up_rx_rdata_11,
  output          up_rx_ready_11,
  output          up_tx_pll_locked_11,
  input           up_tx_rst_11,
  input           up_tx_user_ready_11,
  output          up_tx_rst_done_11,
  input           up_tx_lpm_dfe_n_11,
  input   [ 2:0]  up_tx_rate_11,
  input   [ 1:0]  up_tx_sys_clk_sel_11,
  input   [ 2:0]  up_tx_out_clk_sel_11,
  input   [ 7:0]  up_tx_sel_11,
  input           up_tx_enb_11,
  input   [11:0]  up_tx_addr_11,
  input           up_tx_wr_11,
  input   [15:0]  up_tx_wdata_11,
  output  [15:0]  up_tx_rdata_11,
  output          up_tx_ready_11,

  input           qpll_ref_clk_12,
  input           up_qpll_rst_12,
  input           cpll_ref_clk_12,
  input           up_cpll_rst_12,

  input           rx_12_p,
  input           rx_12_n,
  output          rx_out_clk_12,
  input           rx_clk_12,
  output  [ 3:0]  rx_charisk_12,
  output  [ 3:0]  rx_disperr_12,
  output  [ 3:0]  rx_notintable_12,
  output  [31:0]  rx_data_12,
  input           rx_calign_12,

  output          tx_12_p,
  output          tx_12_n,
  output          tx_out_clk_12,
  input           tx_clk_12,
  input   [ 3:0]  tx_charisk_12,
  input   [31:0]  tx_data_12,

  input   [ 7:0]  up_cm_sel_12,
  input           up_cm_enb_12,
  input   [11:0]  up_cm_addr_12,
  input           up_cm_wr_12,
  input   [15:0]  up_cm_wdata_12,
  output  [15:0]  up_cm_rdata_12,
  output          up_cm_ready_12,
  input   [ 7:0]  up_es_sel_12,
  input           up_es_enb_12,
  input   [11:0]  up_es_addr_12,
  input           up_es_wr_12,
  input   [15:0]  up_es_wdata_12,
  output  [15:0]  up_es_rdata_12,
  output          up_es_ready_12,
  output          up_rx_pll_locked_12,
  input           up_rx_rst_12,
  input           up_rx_user_ready_12,
  output          up_rx_rst_done_12,
  input           up_rx_lpm_dfe_n_12,
  input   [ 2:0]  up_rx_rate_12,
  input   [ 1:0]  up_rx_sys_clk_sel_12,
  input   [ 2:0]  up_rx_out_clk_sel_12,
  input   [ 7:0]  up_rx_sel_12,
  input           up_rx_enb_12,
  input   [11:0]  up_rx_addr_12,
  input           up_rx_wr_12,
  input   [15:0]  up_rx_wdata_12,
  output  [15:0]  up_rx_rdata_12,
  output          up_rx_ready_12,
  output          up_tx_pll_locked_12,
  input           up_tx_rst_12,
  input           up_tx_user_ready_12,
  output          up_tx_rst_done_12,
  input           up_tx_lpm_dfe_n_12,
  input   [ 2:0]  up_tx_rate_12,
  input   [ 1:0]  up_tx_sys_clk_sel_12,
  input   [ 2:0]  up_tx_out_clk_sel_12,
  input   [ 7:0]  up_tx_sel_12,
  input           up_tx_enb_12,
  input   [11:0]  up_tx_addr_12,
  input           up_tx_wr_12,
  input   [15:0]  up_tx_wdata_12,
  output  [15:0]  up_tx_rdata_12,
  output          up_tx_ready_12,

  input           cpll_ref_clk_13,
  input           up_cpll_rst_13,

  input           rx_13_p,
  input           rx_13_n,
  output          rx_out_clk_13,
  input           rx_clk_13,
  output  [ 3:0]  rx_charisk_13,
  output  [ 3:0]  rx_disperr_13,
  output  [ 3:0]  rx_notintable_13,
  output  [31:0]  rx_data_13,
  input           rx_calign_13,

  output          tx_13_p,
  output          tx_13_n,
  output          tx_out_clk_13,
  input           tx_clk_13,
  input   [ 3:0]  tx_charisk_13,
  input   [31:0]  tx_data_13,

  input   [ 7:0]  up_es_sel_13,
  input           up_es_enb_13,
  input   [11:0]  up_es_addr_13,
  input           up_es_wr_13,
  input   [15:0]  up_es_wdata_13,
  output  [15:0]  up_es_rdata_13,
  output          up_es_ready_13,
  output          up_rx_pll_locked_13,
  input           up_rx_rst_13,
  input           up_rx_user_ready_13,
  output          up_rx_rst_done_13,
  input           up_rx_lpm_dfe_n_13,
  input   [ 2:0]  up_rx_rate_13,
  input   [ 1:0]  up_rx_sys_clk_sel_13,
  input   [ 2:0]  up_rx_out_clk_sel_13,
  input   [ 7:0]  up_rx_sel_13,
  input           up_rx_enb_13,
  input   [11:0]  up_rx_addr_13,
  input           up_rx_wr_13,
  input   [15:0]  up_rx_wdata_13,
  output  [15:0]  up_rx_rdata_13,
  output          up_rx_ready_13,
  output          up_tx_pll_locked_13,
  input           up_tx_rst_13,
  input           up_tx_user_ready_13,
  output          up_tx_rst_done_13,
  input           up_tx_lpm_dfe_n_13,
  input   [ 2:0]  up_tx_rate_13,
  input   [ 1:0]  up_tx_sys_clk_sel_13,
  input   [ 2:0]  up_tx_out_clk_sel_13,
  input   [ 7:0]  up_tx_sel_13,
  input           up_tx_enb_13,
  input   [11:0]  up_tx_addr_13,
  input           up_tx_wr_13,
  input   [15:0]  up_tx_wdata_13,
  output  [15:0]  up_tx_rdata_13,
  output          up_tx_ready_13,

  input           cpll_ref_clk_14,
  input           up_cpll_rst_14,

  input           rx_14_p,
  input           rx_14_n,
  output          rx_out_clk_14,
  input           rx_clk_14,
  output  [ 3:0]  rx_charisk_14,
  output  [ 3:0]  rx_disperr_14,
  output  [ 3:0]  rx_notintable_14,
  output  [31:0]  rx_data_14,
  input           rx_calign_14,

  output          tx_14_p,
  output          tx_14_n,
  output          tx_out_clk_14,
  input           tx_clk_14,
  input   [ 3:0]  tx_charisk_14,
  input   [31:0]  tx_data_14,

  input   [ 7:0]  up_es_sel_14,
  input           up_es_enb_14,
  input   [11:0]  up_es_addr_14,
  input           up_es_wr_14,
  input   [15:0]  up_es_wdata_14,
  output  [15:0]  up_es_rdata_14,
  output          up_es_ready_14,
  output          up_rx_pll_locked_14,
  input           up_rx_rst_14,
  input           up_rx_user_ready_14,
  output          up_rx_rst_done_14,
  input           up_rx_lpm_dfe_n_14,
  input   [ 2:0]  up_rx_rate_14,
  input   [ 1:0]  up_rx_sys_clk_sel_14,
  input   [ 2:0]  up_rx_out_clk_sel_14,
  input   [ 7:0]  up_rx_sel_14,
  input           up_rx_enb_14,
  input   [11:0]  up_rx_addr_14,
  input           up_rx_wr_14,
  input   [15:0]  up_rx_wdata_14,
  output  [15:0]  up_rx_rdata_14,
  output          up_rx_ready_14,
  output          up_tx_pll_locked_14,
  input           up_tx_rst_14,
  input           up_tx_user_ready_14,
  output          up_tx_rst_done_14,
  input           up_tx_lpm_dfe_n_14,
  input   [ 2:0]  up_tx_rate_14,
  input   [ 1:0]  up_tx_sys_clk_sel_14,
  input   [ 2:0]  up_tx_out_clk_sel_14,
  input   [ 7:0]  up_tx_sel_14,
  input           up_tx_enb_14,
  input   [11:0]  up_tx_addr_14,
  input           up_tx_wr_14,
  input   [15:0]  up_tx_wdata_14,
  output  [15:0]  up_tx_rdata_14,
  output          up_tx_ready_14,

  input           cpll_ref_clk_15,
  input           up_cpll_rst_15,

  input           rx_15_p,
  input           rx_15_n,
  output          rx_out_clk_15,
  input           rx_clk_15,
  output  [ 3:0]  rx_charisk_15,
  output  [ 3:0]  rx_disperr_15,
  output  [ 3:0]  rx_notintable_15,
  output  [31:0]  rx_data_15,
  input           rx_calign_15,

  output          tx_15_p,
  output          tx_15_n,
  output          tx_out_clk_15,
  input           tx_clk_15,
  input   [ 3:0]  tx_charisk_15,
  input   [31:0]  tx_data_15,

  input   [ 7:0]  up_es_sel_15,
  input           up_es_enb_15,
  input   [11:0]  up_es_addr_15,
  input           up_es_wr_15,
  input   [15:0]  up_es_wdata_15,
  output  [15:0]  up_es_rdata_15,
  output          up_es_ready_15,
  output          up_rx_pll_locked_15,
  input           up_rx_rst_15,
  input           up_rx_user_ready_15,
  output          up_rx_rst_done_15,
  input           up_rx_lpm_dfe_n_15,
  input   [ 2:0]  up_rx_rate_15,
  input   [ 1:0]  up_rx_sys_clk_sel_15,
  input   [ 2:0]  up_rx_out_clk_sel_15,
  input   [ 7:0]  up_rx_sel_15,
  input           up_rx_enb_15,
  input   [11:0]  up_rx_addr_15,
  input           up_rx_wr_15,
  input   [15:0]  up_rx_wdata_15,
  output  [15:0]  up_rx_rdata_15,
  output          up_rx_ready_15,
  output          up_tx_pll_locked_15,
  input           up_tx_rst_15,
  input           up_tx_user_ready_15,
  output          up_tx_rst_done_15,
  input           up_tx_lpm_dfe_n_15,
  input   [ 2:0]  up_tx_rate_15,
  input   [ 1:0]  up_tx_sys_clk_sel_15,
  input   [ 2:0]  up_tx_out_clk_sel_15,
  input   [ 7:0]  up_tx_sel_15,
  input           up_tx_enb_15,
  input   [11:0]  up_tx_addr_15,
  input           up_tx_wr_15,
  input   [15:0]  up_tx_wdata_15,
  output  [15:0]  up_tx_rdata_15,
  output          up_tx_ready_15);

  // parameters

  localparam  integer NUM_OF_LANES = (TX_NUM_OF_LANES > RX_NUM_OF_LANES) ?
    TX_NUM_OF_LANES : RX_NUM_OF_LANES;

  // internal signals

  wire            qpll2ch_clk_0;
  wire            qpll2ch_ref_clk_0;
  wire            qpll2ch_locked_0;
  wire            qpll2ch_clk_4;
  wire            qpll2ch_ref_clk_4;
  wire            qpll2ch_locked_4;
  wire            qpll2ch_clk_8;
  wire            qpll2ch_ref_clk_8;
  wire            qpll2ch_locked_8;
  wire            qpll2ch_clk_12;
  wire            qpll2ch_ref_clk_12;
  wire            qpll2ch_locked_12;

  // instantiations

  generate
  if (NUM_OF_LANES >= 1) begin
  util_adxcvr_xcm #(
    .XCVR_ID (0),
    .XCVR_TYPE (XCVR_TYPE),
    .QPLL_REFCLK_DIV (QPLL_REFCLK_DIV),
    .QPLL_FBDIV_RATIO (QPLL_FBDIV_RATIO),
    .QPLL_CFG (QPLL_CFG),
    .QPLL_FBDIV (QPLL_FBDIV))
  i_xcm_0 (
    .qpll_ref_clk (qpll_ref_clk_0),
    .qpll2ch_clk (qpll2ch_clk_0),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_0),
    .qpll2ch_locked (qpll2ch_locked_0),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_qpll_rst (up_qpll_rst_0),
    .up_cm_sel (up_cm_sel_0),
    .up_cm_enb (up_cm_enb_0),
    .up_cm_addr (up_cm_addr_0),
    .up_cm_wr (up_cm_wr_0),
    .up_cm_wdata (up_cm_wdata_0),
    .up_cm_rdata (up_cm_rdata_0),
    .up_cm_ready (up_cm_ready_0));
  end else begin
  assign qpll2ch_clk_0 = 1'd0;
  assign qpll2ch_ref_clk_0 = 1'd0;
  assign qpll2ch_locked_0 = 1'd0;
  assign up_cm_rdata_0 = 16'd0;
  assign up_cm_ready_0 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 1) begin
  util_adxcvr_xch #(
    .XCVR_ID (0),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_0 (
    .qpll2ch_clk (qpll2ch_clk_0),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_0),
    .qpll2ch_locked (qpll2ch_locked_0),
    .cpll_ref_clk (cpll_ref_clk_0),
    .up_cpll_rst (up_cpll_rst_0),
    .rx_p (rx_0_p),
    .rx_n (rx_0_n),
    .rx_out_clk (rx_out_clk_0),
    .rx_clk (rx_clk_0),
    .rx_charisk (rx_charisk_0),
    .rx_disperr (rx_disperr_0),
    .rx_notintable (rx_notintable_0),
    .rx_data (rx_data_0),
    .rx_calign (rx_calign_0),
    .tx_p (tx_0_p),
    .tx_n (tx_0_n),
    .tx_out_clk (tx_out_clk_0),
    .tx_clk (tx_clk_0),
    .tx_charisk (tx_charisk_0),
    .tx_data (tx_data_0),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_0),
    .up_es_enb (up_es_enb_0),
    .up_es_addr (up_es_addr_0),
    .up_es_wr (up_es_wr_0),
    .up_es_wdata (up_es_wdata_0),
    .up_es_rdata (up_es_rdata_0),
    .up_es_ready (up_es_ready_0),
    .up_rx_pll_locked (up_rx_pll_locked_0),
    .up_rx_rst (up_rx_rst_0),
    .up_rx_user_ready (up_rx_user_ready_0),
    .up_rx_rst_done (up_rx_rst_done_0),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_0),
    .up_rx_rate (up_rx_rate_0),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_0),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_0),
    .up_rx_sel (up_rx_sel_0),
    .up_rx_enb (up_rx_enb_0),
    .up_rx_addr (up_rx_addr_0),
    .up_rx_wr (up_rx_wr_0),
    .up_rx_wdata (up_rx_wdata_0),
    .up_rx_rdata (up_rx_rdata_0),
    .up_rx_ready (up_rx_ready_0),
    .up_tx_pll_locked (up_tx_pll_locked_0),
    .up_tx_rst (up_tx_rst_0),
    .up_tx_user_ready (up_tx_user_ready_0),
    .up_tx_rst_done (up_tx_rst_done_0),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_0),
    .up_tx_rate (up_tx_rate_0),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_0),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_0),
    .up_tx_sel (up_tx_sel_0),
    .up_tx_enb (up_tx_enb_0),
    .up_tx_addr (up_tx_addr_0),
    .up_tx_wr (up_tx_wr_0),
    .up_tx_wdata (up_tx_wdata_0),
    .up_tx_rdata (up_tx_rdata_0),
    .up_tx_ready (up_tx_ready_0));
  end else begin
  assign rx_out_clk_0 = 1'd0;
  assign rx_charisk_0 = 4'd0;
  assign rx_disperr_0 = 4'd0;
  assign rx_notintable_0 = 4'd0;
  assign rx_data_0 = 32'd0;
  assign tx_0_p = 1'd0;
  assign tx_0_n = 1'd0;
  assign tx_out_clk_0 = 1'd0;
  assign up_es_rdata_0 = 16'd0;
  assign up_es_ready_0 = 1'd0;
  assign up_rx_pll_locked_0 = 1'd0;
  assign up_rx_rst_done_0 = 1'd0;
  assign up_rx_rdata_0 = 16'd0;
  assign up_rx_ready_0 = 1'd0;
  assign up_tx_pll_locked_0 = 1'd0;
  assign up_tx_rst_done_0 = 1'd0;
  assign up_tx_rdata_0 = 16'd0;
  assign up_tx_ready_0 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 2) begin
  util_adxcvr_xch #(
    .XCVR_ID (1),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_1 (
    .qpll2ch_clk (qpll2ch_clk_0),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_0),
    .qpll2ch_locked (qpll2ch_locked_0),
    .cpll_ref_clk (cpll_ref_clk_1),
    .up_cpll_rst (up_cpll_rst_1),
    .rx_p (rx_1_p),
    .rx_n (rx_1_n),
    .rx_out_clk (rx_out_clk_1),
    .rx_clk (rx_clk_1),
    .rx_charisk (rx_charisk_1),
    .rx_disperr (rx_disperr_1),
    .rx_notintable (rx_notintable_1),
    .rx_data (rx_data_1),
    .rx_calign (rx_calign_1),
    .tx_p (tx_1_p),
    .tx_n (tx_1_n),
    .tx_out_clk (tx_out_clk_1),
    .tx_clk (tx_clk_1),
    .tx_charisk (tx_charisk_1),
    .tx_data (tx_data_1),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_1),
    .up_es_enb (up_es_enb_1),
    .up_es_addr (up_es_addr_1),
    .up_es_wr (up_es_wr_1),
    .up_es_wdata (up_es_wdata_1),
    .up_es_rdata (up_es_rdata_1),
    .up_es_ready (up_es_ready_1),
    .up_rx_pll_locked (up_rx_pll_locked_1),
    .up_rx_rst (up_rx_rst_1),
    .up_rx_user_ready (up_rx_user_ready_1),
    .up_rx_rst_done (up_rx_rst_done_1),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_1),
    .up_rx_rate (up_rx_rate_1),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_1),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_1),
    .up_rx_sel (up_rx_sel_1),
    .up_rx_enb (up_rx_enb_1),
    .up_rx_addr (up_rx_addr_1),
    .up_rx_wr (up_rx_wr_1),
    .up_rx_wdata (up_rx_wdata_1),
    .up_rx_rdata (up_rx_rdata_1),
    .up_rx_ready (up_rx_ready_1),
    .up_tx_pll_locked (up_tx_pll_locked_1),
    .up_tx_rst (up_tx_rst_1),
    .up_tx_user_ready (up_tx_user_ready_1),
    .up_tx_rst_done (up_tx_rst_done_1),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_1),
    .up_tx_rate (up_tx_rate_1),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_1),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_1),
    .up_tx_sel (up_tx_sel_1),
    .up_tx_enb (up_tx_enb_1),
    .up_tx_addr (up_tx_addr_1),
    .up_tx_wr (up_tx_wr_1),
    .up_tx_wdata (up_tx_wdata_1),
    .up_tx_rdata (up_tx_rdata_1),
    .up_tx_ready (up_tx_ready_1));
  end else begin
  assign rx_out_clk_1 = 1'd0;
  assign rx_charisk_1 = 4'd0;
  assign rx_disperr_1 = 4'd0;
  assign rx_notintable_1 = 4'd0;
  assign rx_data_1 = 32'd0;
  assign tx_1_p = 1'd0;
  assign tx_1_n = 1'd0;
  assign tx_out_clk_1 = 1'd0;
  assign up_es_rdata_1 = 16'd0;
  assign up_es_ready_1 = 1'd0;
  assign up_rx_pll_locked_1 = 1'd0;
  assign up_rx_rst_done_1 = 1'd0;
  assign up_rx_rdata_1 = 16'd0;
  assign up_rx_ready_1 = 1'd0;
  assign up_tx_pll_locked_1 = 1'd0;
  assign up_tx_rst_done_1 = 1'd0;
  assign up_tx_rdata_1 = 16'd0;
  assign up_tx_ready_1 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 3) begin
  util_adxcvr_xch #(
    .XCVR_ID (2),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_2 (
    .qpll2ch_clk (qpll2ch_clk_0),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_0),
    .qpll2ch_locked (qpll2ch_locked_0),
    .cpll_ref_clk (cpll_ref_clk_2),
    .up_cpll_rst (up_cpll_rst_2),
    .rx_p (rx_2_p),
    .rx_n (rx_2_n),
    .rx_out_clk (rx_out_clk_2),
    .rx_clk (rx_clk_2),
    .rx_charisk (rx_charisk_2),
    .rx_disperr (rx_disperr_2),
    .rx_notintable (rx_notintable_2),
    .rx_data (rx_data_2),
    .rx_calign (rx_calign_2),
    .tx_p (tx_2_p),
    .tx_n (tx_2_n),
    .tx_out_clk (tx_out_clk_2),
    .tx_clk (tx_clk_2),
    .tx_charisk (tx_charisk_2),
    .tx_data (tx_data_2),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_2),
    .up_es_enb (up_es_enb_2),
    .up_es_addr (up_es_addr_2),
    .up_es_wr (up_es_wr_2),
    .up_es_wdata (up_es_wdata_2),
    .up_es_rdata (up_es_rdata_2),
    .up_es_ready (up_es_ready_2),
    .up_rx_pll_locked (up_rx_pll_locked_2),
    .up_rx_rst (up_rx_rst_2),
    .up_rx_user_ready (up_rx_user_ready_2),
    .up_rx_rst_done (up_rx_rst_done_2),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_2),
    .up_rx_rate (up_rx_rate_2),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_2),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_2),
    .up_rx_sel (up_rx_sel_2),
    .up_rx_enb (up_rx_enb_2),
    .up_rx_addr (up_rx_addr_2),
    .up_rx_wr (up_rx_wr_2),
    .up_rx_wdata (up_rx_wdata_2),
    .up_rx_rdata (up_rx_rdata_2),
    .up_rx_ready (up_rx_ready_2),
    .up_tx_pll_locked (up_tx_pll_locked_2),
    .up_tx_rst (up_tx_rst_2),
    .up_tx_user_ready (up_tx_user_ready_2),
    .up_tx_rst_done (up_tx_rst_done_2),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_2),
    .up_tx_rate (up_tx_rate_2),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_2),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_2),
    .up_tx_sel (up_tx_sel_2),
    .up_tx_enb (up_tx_enb_2),
    .up_tx_addr (up_tx_addr_2),
    .up_tx_wr (up_tx_wr_2),
    .up_tx_wdata (up_tx_wdata_2),
    .up_tx_rdata (up_tx_rdata_2),
    .up_tx_ready (up_tx_ready_2));
  end else begin
  assign rx_out_clk_2 = 1'd0;
  assign rx_charisk_2 = 4'd0;
  assign rx_disperr_2 = 4'd0;
  assign rx_notintable_2 = 4'd0;
  assign rx_data_2 = 32'd0;
  assign tx_2_p = 1'd0;
  assign tx_2_n = 1'd0;
  assign tx_out_clk_2 = 1'd0;
  assign up_es_rdata_2 = 16'd0;
  assign up_es_ready_2 = 1'd0;
  assign up_rx_pll_locked_2 = 1'd0;
  assign up_rx_rst_done_2 = 1'd0;
  assign up_rx_rdata_2 = 16'd0;
  assign up_rx_ready_2 = 1'd0;
  assign up_tx_pll_locked_2 = 1'd0;
  assign up_tx_rst_done_2 = 1'd0;
  assign up_tx_rdata_2 = 16'd0;
  assign up_tx_ready_2 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 4) begin
  util_adxcvr_xch #(
    .XCVR_ID (3),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_3 (
    .qpll2ch_clk (qpll2ch_clk_0),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_0),
    .qpll2ch_locked (qpll2ch_locked_0),
    .cpll_ref_clk (cpll_ref_clk_3),
    .up_cpll_rst (up_cpll_rst_3),
    .rx_p (rx_3_p),
    .rx_n (rx_3_n),
    .rx_out_clk (rx_out_clk_3),
    .rx_clk (rx_clk_3),
    .rx_charisk (rx_charisk_3),
    .rx_disperr (rx_disperr_3),
    .rx_notintable (rx_notintable_3),
    .rx_data (rx_data_3),
    .rx_calign (rx_calign_3),
    .tx_p (tx_3_p),
    .tx_n (tx_3_n),
    .tx_out_clk (tx_out_clk_3),
    .tx_clk (tx_clk_3),
    .tx_charisk (tx_charisk_3),
    .tx_data (tx_data_3),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_3),
    .up_es_enb (up_es_enb_3),
    .up_es_addr (up_es_addr_3),
    .up_es_wr (up_es_wr_3),
    .up_es_wdata (up_es_wdata_3),
    .up_es_rdata (up_es_rdata_3),
    .up_es_ready (up_es_ready_3),
    .up_rx_pll_locked (up_rx_pll_locked_3),
    .up_rx_rst (up_rx_rst_3),
    .up_rx_user_ready (up_rx_user_ready_3),
    .up_rx_rst_done (up_rx_rst_done_3),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_3),
    .up_rx_rate (up_rx_rate_3),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_3),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_3),
    .up_rx_sel (up_rx_sel_3),
    .up_rx_enb (up_rx_enb_3),
    .up_rx_addr (up_rx_addr_3),
    .up_rx_wr (up_rx_wr_3),
    .up_rx_wdata (up_rx_wdata_3),
    .up_rx_rdata (up_rx_rdata_3),
    .up_rx_ready (up_rx_ready_3),
    .up_tx_pll_locked (up_tx_pll_locked_3),
    .up_tx_rst (up_tx_rst_3),
    .up_tx_user_ready (up_tx_user_ready_3),
    .up_tx_rst_done (up_tx_rst_done_3),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_3),
    .up_tx_rate (up_tx_rate_3),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_3),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_3),
    .up_tx_sel (up_tx_sel_3),
    .up_tx_enb (up_tx_enb_3),
    .up_tx_addr (up_tx_addr_3),
    .up_tx_wr (up_tx_wr_3),
    .up_tx_wdata (up_tx_wdata_3),
    .up_tx_rdata (up_tx_rdata_3),
    .up_tx_ready (up_tx_ready_3));
  end else begin
  assign rx_out_clk_3 = 1'd0;
  assign rx_charisk_3 = 4'd0;
  assign rx_disperr_3 = 4'd0;
  assign rx_notintable_3 = 4'd0;
  assign rx_data_3 = 32'd0;
  assign tx_3_p = 1'd0;
  assign tx_3_n = 1'd0;
  assign tx_out_clk_3 = 1'd0;
  assign up_es_rdata_3 = 16'd0;
  assign up_es_ready_3 = 1'd0;
  assign up_rx_pll_locked_3 = 1'd0;
  assign up_rx_rst_done_3 = 1'd0;
  assign up_rx_rdata_3 = 16'd0;
  assign up_rx_ready_3 = 1'd0;
  assign up_tx_pll_locked_3 = 1'd0;
  assign up_tx_rst_done_3 = 1'd0;
  assign up_tx_rdata_3 = 16'd0;
  assign up_tx_ready_3 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 5) begin
  util_adxcvr_xcm #(
    .XCVR_ID (4),
    .XCVR_TYPE (XCVR_TYPE),
    .QPLL_REFCLK_DIV (QPLL_REFCLK_DIV),
    .QPLL_FBDIV_RATIO (QPLL_FBDIV_RATIO),
    .QPLL_CFG (QPLL_CFG),
    .QPLL_FBDIV (QPLL_FBDIV))
  i_xcm_4 (
    .qpll_ref_clk (qpll_ref_clk_4),
    .qpll2ch_clk (qpll2ch_clk_4),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_4),
    .qpll2ch_locked (qpll2ch_locked_4),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_qpll_rst (up_qpll_rst_4),
    .up_cm_sel (up_cm_sel_4),
    .up_cm_enb (up_cm_enb_4),
    .up_cm_addr (up_cm_addr_4),
    .up_cm_wr (up_cm_wr_4),
    .up_cm_wdata (up_cm_wdata_4),
    .up_cm_rdata (up_cm_rdata_4),
    .up_cm_ready (up_cm_ready_4));
  end else begin
  assign qpll2ch_clk_4 = 1'd0;
  assign qpll2ch_ref_clk_4 = 1'd0;
  assign qpll2ch_locked_4 = 1'd0;
  assign up_cm_rdata_4 = 16'd0;
  assign up_cm_ready_4 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 5) begin
  util_adxcvr_xch #(
    .XCVR_ID (4),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_4 (
    .qpll2ch_clk (qpll2ch_clk_4),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_4),
    .qpll2ch_locked (qpll2ch_locked_4),
    .cpll_ref_clk (cpll_ref_clk_4),
    .up_cpll_rst (up_cpll_rst_4),
    .rx_p (rx_4_p),
    .rx_n (rx_4_n),
    .rx_out_clk (rx_out_clk_4),
    .rx_clk (rx_clk_4),
    .rx_charisk (rx_charisk_4),
    .rx_disperr (rx_disperr_4),
    .rx_notintable (rx_notintable_4),
    .rx_data (rx_data_4),
    .rx_calign (rx_calign_4),
    .tx_p (tx_4_p),
    .tx_n (tx_4_n),
    .tx_out_clk (tx_out_clk_4),
    .tx_clk (tx_clk_4),
    .tx_charisk (tx_charisk_4),
    .tx_data (tx_data_4),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_4),
    .up_es_enb (up_es_enb_4),
    .up_es_addr (up_es_addr_4),
    .up_es_wr (up_es_wr_4),
    .up_es_wdata (up_es_wdata_4),
    .up_es_rdata (up_es_rdata_4),
    .up_es_ready (up_es_ready_4),
    .up_rx_pll_locked (up_rx_pll_locked_4),
    .up_rx_rst (up_rx_rst_4),
    .up_rx_user_ready (up_rx_user_ready_4),
    .up_rx_rst_done (up_rx_rst_done_4),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_4),
    .up_rx_rate (up_rx_rate_4),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_4),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_4),
    .up_rx_sel (up_rx_sel_4),
    .up_rx_enb (up_rx_enb_4),
    .up_rx_addr (up_rx_addr_4),
    .up_rx_wr (up_rx_wr_4),
    .up_rx_wdata (up_rx_wdata_4),
    .up_rx_rdata (up_rx_rdata_4),
    .up_rx_ready (up_rx_ready_4),
    .up_tx_pll_locked (up_tx_pll_locked_4),
    .up_tx_rst (up_tx_rst_4),
    .up_tx_user_ready (up_tx_user_ready_4),
    .up_tx_rst_done (up_tx_rst_done_4),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_4),
    .up_tx_rate (up_tx_rate_4),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_4),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_4),
    .up_tx_sel (up_tx_sel_4),
    .up_tx_enb (up_tx_enb_4),
    .up_tx_addr (up_tx_addr_4),
    .up_tx_wr (up_tx_wr_4),
    .up_tx_wdata (up_tx_wdata_4),
    .up_tx_rdata (up_tx_rdata_4),
    .up_tx_ready (up_tx_ready_4));
  end else begin
  assign rx_out_clk_4 = 1'd0;
  assign rx_charisk_4 = 4'd0;
  assign rx_disperr_4 = 4'd0;
  assign rx_notintable_4 = 4'd0;
  assign rx_data_4 = 32'd0;
  assign tx_4_p = 1'd0;
  assign tx_4_n = 1'd0;
  assign tx_out_clk_4 = 1'd0;
  assign up_es_rdata_4 = 16'd0;
  assign up_es_ready_4 = 1'd0;
  assign up_rx_pll_locked_4 = 1'd0;
  assign up_rx_rst_done_4 = 1'd0;
  assign up_rx_rdata_4 = 16'd0;
  assign up_rx_ready_4 = 1'd0;
  assign up_tx_pll_locked_4 = 1'd0;
  assign up_tx_rst_done_4 = 1'd0;
  assign up_tx_rdata_4 = 16'd0;
  assign up_tx_ready_4 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 6) begin
  util_adxcvr_xch #(
    .XCVR_ID (5),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_5 (
    .qpll2ch_clk (qpll2ch_clk_4),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_4),
    .qpll2ch_locked (qpll2ch_locked_4),
    .cpll_ref_clk (cpll_ref_clk_5),
    .up_cpll_rst (up_cpll_rst_5),
    .rx_p (rx_5_p),
    .rx_n (rx_5_n),
    .rx_out_clk (rx_out_clk_5),
    .rx_clk (rx_clk_5),
    .rx_charisk (rx_charisk_5),
    .rx_disperr (rx_disperr_5),
    .rx_notintable (rx_notintable_5),
    .rx_data (rx_data_5),
    .rx_calign (rx_calign_5),
    .tx_p (tx_5_p),
    .tx_n (tx_5_n),
    .tx_out_clk (tx_out_clk_5),
    .tx_clk (tx_clk_5),
    .tx_charisk (tx_charisk_5),
    .tx_data (tx_data_5),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_5),
    .up_es_enb (up_es_enb_5),
    .up_es_addr (up_es_addr_5),
    .up_es_wr (up_es_wr_5),
    .up_es_wdata (up_es_wdata_5),
    .up_es_rdata (up_es_rdata_5),
    .up_es_ready (up_es_ready_5),
    .up_rx_pll_locked (up_rx_pll_locked_5),
    .up_rx_rst (up_rx_rst_5),
    .up_rx_user_ready (up_rx_user_ready_5),
    .up_rx_rst_done (up_rx_rst_done_5),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_5),
    .up_rx_rate (up_rx_rate_5),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_5),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_5),
    .up_rx_sel (up_rx_sel_5),
    .up_rx_enb (up_rx_enb_5),
    .up_rx_addr (up_rx_addr_5),
    .up_rx_wr (up_rx_wr_5),
    .up_rx_wdata (up_rx_wdata_5),
    .up_rx_rdata (up_rx_rdata_5),
    .up_rx_ready (up_rx_ready_5),
    .up_tx_pll_locked (up_tx_pll_locked_5),
    .up_tx_rst (up_tx_rst_5),
    .up_tx_user_ready (up_tx_user_ready_5),
    .up_tx_rst_done (up_tx_rst_done_5),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_5),
    .up_tx_rate (up_tx_rate_5),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_5),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_5),
    .up_tx_sel (up_tx_sel_5),
    .up_tx_enb (up_tx_enb_5),
    .up_tx_addr (up_tx_addr_5),
    .up_tx_wr (up_tx_wr_5),
    .up_tx_wdata (up_tx_wdata_5),
    .up_tx_rdata (up_tx_rdata_5),
    .up_tx_ready (up_tx_ready_5));
  end else begin
  assign rx_out_clk_5 = 1'd0;
  assign rx_charisk_5 = 4'd0;
  assign rx_disperr_5 = 4'd0;
  assign rx_notintable_5 = 4'd0;
  assign rx_data_5 = 32'd0;
  assign tx_5_p = 1'd0;
  assign tx_5_n = 1'd0;
  assign tx_out_clk_5 = 1'd0;
  assign up_es_rdata_5 = 16'd0;
  assign up_es_ready_5 = 1'd0;
  assign up_rx_pll_locked_5 = 1'd0;
  assign up_rx_rst_done_5 = 1'd0;
  assign up_rx_rdata_5 = 16'd0;
  assign up_rx_ready_5 = 1'd0;
  assign up_tx_pll_locked_5 = 1'd0;
  assign up_tx_rst_done_5 = 1'd0;
  assign up_tx_rdata_5 = 16'd0;
  assign up_tx_ready_5 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 7) begin
  util_adxcvr_xch #(
    .XCVR_ID (6),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_6 (
    .qpll2ch_clk (qpll2ch_clk_4),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_4),
    .qpll2ch_locked (qpll2ch_locked_4),
    .cpll_ref_clk (cpll_ref_clk_6),
    .up_cpll_rst (up_cpll_rst_6),
    .rx_p (rx_6_p),
    .rx_n (rx_6_n),
    .rx_out_clk (rx_out_clk_6),
    .rx_clk (rx_clk_6),
    .rx_charisk (rx_charisk_6),
    .rx_disperr (rx_disperr_6),
    .rx_notintable (rx_notintable_6),
    .rx_data (rx_data_6),
    .rx_calign (rx_calign_6),
    .tx_p (tx_6_p),
    .tx_n (tx_6_n),
    .tx_out_clk (tx_out_clk_6),
    .tx_clk (tx_clk_6),
    .tx_charisk (tx_charisk_6),
    .tx_data (tx_data_6),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_6),
    .up_es_enb (up_es_enb_6),
    .up_es_addr (up_es_addr_6),
    .up_es_wr (up_es_wr_6),
    .up_es_wdata (up_es_wdata_6),
    .up_es_rdata (up_es_rdata_6),
    .up_es_ready (up_es_ready_6),
    .up_rx_pll_locked (up_rx_pll_locked_6),
    .up_rx_rst (up_rx_rst_6),
    .up_rx_user_ready (up_rx_user_ready_6),
    .up_rx_rst_done (up_rx_rst_done_6),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_6),
    .up_rx_rate (up_rx_rate_6),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_6),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_6),
    .up_rx_sel (up_rx_sel_6),
    .up_rx_enb (up_rx_enb_6),
    .up_rx_addr (up_rx_addr_6),
    .up_rx_wr (up_rx_wr_6),
    .up_rx_wdata (up_rx_wdata_6),
    .up_rx_rdata (up_rx_rdata_6),
    .up_rx_ready (up_rx_ready_6),
    .up_tx_pll_locked (up_tx_pll_locked_6),
    .up_tx_rst (up_tx_rst_6),
    .up_tx_user_ready (up_tx_user_ready_6),
    .up_tx_rst_done (up_tx_rst_done_6),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_6),
    .up_tx_rate (up_tx_rate_6),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_6),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_6),
    .up_tx_sel (up_tx_sel_6),
    .up_tx_enb (up_tx_enb_6),
    .up_tx_addr (up_tx_addr_6),
    .up_tx_wr (up_tx_wr_6),
    .up_tx_wdata (up_tx_wdata_6),
    .up_tx_rdata (up_tx_rdata_6),
    .up_tx_ready (up_tx_ready_6));
  end else begin
  assign rx_out_clk_6 = 1'd0;
  assign rx_charisk_6 = 4'd0;
  assign rx_disperr_6 = 4'd0;
  assign rx_notintable_6 = 4'd0;
  assign rx_data_6 = 32'd0;
  assign tx_6_p = 1'd0;
  assign tx_6_n = 1'd0;
  assign tx_out_clk_6 = 1'd0;
  assign up_es_rdata_6 = 16'd0;
  assign up_es_ready_6 = 1'd0;
  assign up_rx_pll_locked_6 = 1'd0;
  assign up_rx_rst_done_6 = 1'd0;
  assign up_rx_rdata_6 = 16'd0;
  assign up_rx_ready_6 = 1'd0;
  assign up_tx_pll_locked_6 = 1'd0;
  assign up_tx_rst_done_6 = 1'd0;
  assign up_tx_rdata_6 = 16'd0;
  assign up_tx_ready_6 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 8) begin
  util_adxcvr_xch #(
    .XCVR_ID (7),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_7 (
    .qpll2ch_clk (qpll2ch_clk_4),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_4),
    .qpll2ch_locked (qpll2ch_locked_4),
    .cpll_ref_clk (cpll_ref_clk_7),
    .up_cpll_rst (up_cpll_rst_7),
    .rx_p (rx_7_p),
    .rx_n (rx_7_n),
    .rx_out_clk (rx_out_clk_7),
    .rx_clk (rx_clk_7),
    .rx_charisk (rx_charisk_7),
    .rx_disperr (rx_disperr_7),
    .rx_notintable (rx_notintable_7),
    .rx_data (rx_data_7),
    .rx_calign (rx_calign_7),
    .tx_p (tx_7_p),
    .tx_n (tx_7_n),
    .tx_out_clk (tx_out_clk_7),
    .tx_clk (tx_clk_7),
    .tx_charisk (tx_charisk_7),
    .tx_data (tx_data_7),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_7),
    .up_es_enb (up_es_enb_7),
    .up_es_addr (up_es_addr_7),
    .up_es_wr (up_es_wr_7),
    .up_es_wdata (up_es_wdata_7),
    .up_es_rdata (up_es_rdata_7),
    .up_es_ready (up_es_ready_7),
    .up_rx_pll_locked (up_rx_pll_locked_7),
    .up_rx_rst (up_rx_rst_7),
    .up_rx_user_ready (up_rx_user_ready_7),
    .up_rx_rst_done (up_rx_rst_done_7),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_7),
    .up_rx_rate (up_rx_rate_7),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_7),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_7),
    .up_rx_sel (up_rx_sel_7),
    .up_rx_enb (up_rx_enb_7),
    .up_rx_addr (up_rx_addr_7),
    .up_rx_wr (up_rx_wr_7),
    .up_rx_wdata (up_rx_wdata_7),
    .up_rx_rdata (up_rx_rdata_7),
    .up_rx_ready (up_rx_ready_7),
    .up_tx_pll_locked (up_tx_pll_locked_7),
    .up_tx_rst (up_tx_rst_7),
    .up_tx_user_ready (up_tx_user_ready_7),
    .up_tx_rst_done (up_tx_rst_done_7),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_7),
    .up_tx_rate (up_tx_rate_7),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_7),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_7),
    .up_tx_sel (up_tx_sel_7),
    .up_tx_enb (up_tx_enb_7),
    .up_tx_addr (up_tx_addr_7),
    .up_tx_wr (up_tx_wr_7),
    .up_tx_wdata (up_tx_wdata_7),
    .up_tx_rdata (up_tx_rdata_7),
    .up_tx_ready (up_tx_ready_7));
  end else begin
  assign rx_out_clk_7 = 1'd0;
  assign rx_charisk_7 = 4'd0;
  assign rx_disperr_7 = 4'd0;
  assign rx_notintable_7 = 4'd0;
  assign rx_data_7 = 32'd0;
  assign tx_7_p = 1'd0;
  assign tx_7_n = 1'd0;
  assign tx_out_clk_7 = 1'd0;
  assign up_es_rdata_7 = 16'd0;
  assign up_es_ready_7 = 1'd0;
  assign up_rx_pll_locked_7 = 1'd0;
  assign up_rx_rst_done_7 = 1'd0;
  assign up_rx_rdata_7 = 16'd0;
  assign up_rx_ready_7 = 1'd0;
  assign up_tx_pll_locked_7 = 1'd0;
  assign up_tx_rst_done_7 = 1'd0;
  assign up_tx_rdata_7 = 16'd0;
  assign up_tx_ready_7 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 9) begin
  util_adxcvr_xcm #(
    .XCVR_ID (8),
    .XCVR_TYPE (XCVR_TYPE),
    .QPLL_REFCLK_DIV (QPLL_REFCLK_DIV),
    .QPLL_FBDIV_RATIO (QPLL_FBDIV_RATIO),
    .QPLL_CFG (QPLL_CFG),
    .QPLL_FBDIV (QPLL_FBDIV))
  i_xcm_8 (
    .qpll_ref_clk (qpll_ref_clk_8),
    .qpll2ch_clk (qpll2ch_clk_8),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_8),
    .qpll2ch_locked (qpll2ch_locked_8),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_qpll_rst (up_qpll_rst_8),
    .up_cm_sel (up_cm_sel_8),
    .up_cm_enb (up_cm_enb_8),
    .up_cm_addr (up_cm_addr_8),
    .up_cm_wr (up_cm_wr_8),
    .up_cm_wdata (up_cm_wdata_8),
    .up_cm_rdata (up_cm_rdata_8),
    .up_cm_ready (up_cm_ready_8));
  end else begin
  assign qpll2ch_clk_8 = 1'd0;
  assign qpll2ch_ref_clk_8 = 1'd0;
  assign qpll2ch_locked_8 = 1'd0;
  assign up_cm_rdata_8 = 16'd0;
  assign up_cm_ready_8 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 9) begin
  util_adxcvr_xch #(
    .XCVR_ID (8),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_8 (
    .qpll2ch_clk (qpll2ch_clk_8),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_8),
    .qpll2ch_locked (qpll2ch_locked_8),
    .cpll_ref_clk (cpll_ref_clk_8),
    .up_cpll_rst (up_cpll_rst_8),
    .rx_p (rx_8_p),
    .rx_n (rx_8_n),
    .rx_out_clk (rx_out_clk_8),
    .rx_clk (rx_clk_8),
    .rx_charisk (rx_charisk_8),
    .rx_disperr (rx_disperr_8),
    .rx_notintable (rx_notintable_8),
    .rx_data (rx_data_8),
    .rx_calign (rx_calign_8),
    .tx_p (tx_8_p),
    .tx_n (tx_8_n),
    .tx_out_clk (tx_out_clk_8),
    .tx_clk (tx_clk_8),
    .tx_charisk (tx_charisk_8),
    .tx_data (tx_data_8),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_8),
    .up_es_enb (up_es_enb_8),
    .up_es_addr (up_es_addr_8),
    .up_es_wr (up_es_wr_8),
    .up_es_wdata (up_es_wdata_8),
    .up_es_rdata (up_es_rdata_8),
    .up_es_ready (up_es_ready_8),
    .up_rx_pll_locked (up_rx_pll_locked_8),
    .up_rx_rst (up_rx_rst_8),
    .up_rx_user_ready (up_rx_user_ready_8),
    .up_rx_rst_done (up_rx_rst_done_8),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_8),
    .up_rx_rate (up_rx_rate_8),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_8),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_8),
    .up_rx_sel (up_rx_sel_8),
    .up_rx_enb (up_rx_enb_8),
    .up_rx_addr (up_rx_addr_8),
    .up_rx_wr (up_rx_wr_8),
    .up_rx_wdata (up_rx_wdata_8),
    .up_rx_rdata (up_rx_rdata_8),
    .up_rx_ready (up_rx_ready_8),
    .up_tx_pll_locked (up_tx_pll_locked_8),
    .up_tx_rst (up_tx_rst_8),
    .up_tx_user_ready (up_tx_user_ready_8),
    .up_tx_rst_done (up_tx_rst_done_8),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_8),
    .up_tx_rate (up_tx_rate_8),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_8),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_8),
    .up_tx_sel (up_tx_sel_8),
    .up_tx_enb (up_tx_enb_8),
    .up_tx_addr (up_tx_addr_8),
    .up_tx_wr (up_tx_wr_8),
    .up_tx_wdata (up_tx_wdata_8),
    .up_tx_rdata (up_tx_rdata_8),
    .up_tx_ready (up_tx_ready_8));
  end else begin
  assign rx_out_clk_8 = 1'd0;
  assign rx_charisk_8 = 4'd0;
  assign rx_disperr_8 = 4'd0;
  assign rx_notintable_8 = 4'd0;
  assign rx_data_8 = 32'd0;
  assign tx_8_p = 1'd0;
  assign tx_8_n = 1'd0;
  assign tx_out_clk_8 = 1'd0;
  assign up_es_rdata_8 = 16'd0;
  assign up_es_ready_8 = 1'd0;
  assign up_rx_pll_locked_8 = 1'd0;
  assign up_rx_rst_done_8 = 1'd0;
  assign up_rx_rdata_8 = 16'd0;
  assign up_rx_ready_8 = 1'd0;
  assign up_tx_pll_locked_8 = 1'd0;
  assign up_tx_rst_done_8 = 1'd0;
  assign up_tx_rdata_8 = 16'd0;
  assign up_tx_ready_8 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 10) begin
  util_adxcvr_xch #(
    .XCVR_ID (9),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_9 (
    .qpll2ch_clk (qpll2ch_clk_8),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_8),
    .qpll2ch_locked (qpll2ch_locked_8),
    .cpll_ref_clk (cpll_ref_clk_9),
    .up_cpll_rst (up_cpll_rst_9),
    .rx_p (rx_9_p),
    .rx_n (rx_9_n),
    .rx_out_clk (rx_out_clk_9),
    .rx_clk (rx_clk_9),
    .rx_charisk (rx_charisk_9),
    .rx_disperr (rx_disperr_9),
    .rx_notintable (rx_notintable_9),
    .rx_data (rx_data_9),
    .rx_calign (rx_calign_9),
    .tx_p (tx_9_p),
    .tx_n (tx_9_n),
    .tx_out_clk (tx_out_clk_9),
    .tx_clk (tx_clk_9),
    .tx_charisk (tx_charisk_9),
    .tx_data (tx_data_9),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_9),
    .up_es_enb (up_es_enb_9),
    .up_es_addr (up_es_addr_9),
    .up_es_wr (up_es_wr_9),
    .up_es_wdata (up_es_wdata_9),
    .up_es_rdata (up_es_rdata_9),
    .up_es_ready (up_es_ready_9),
    .up_rx_pll_locked (up_rx_pll_locked_9),
    .up_rx_rst (up_rx_rst_9),
    .up_rx_user_ready (up_rx_user_ready_9),
    .up_rx_rst_done (up_rx_rst_done_9),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_9),
    .up_rx_rate (up_rx_rate_9),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_9),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_9),
    .up_rx_sel (up_rx_sel_9),
    .up_rx_enb (up_rx_enb_9),
    .up_rx_addr (up_rx_addr_9),
    .up_rx_wr (up_rx_wr_9),
    .up_rx_wdata (up_rx_wdata_9),
    .up_rx_rdata (up_rx_rdata_9),
    .up_rx_ready (up_rx_ready_9),
    .up_tx_pll_locked (up_tx_pll_locked_9),
    .up_tx_rst (up_tx_rst_9),
    .up_tx_user_ready (up_tx_user_ready_9),
    .up_tx_rst_done (up_tx_rst_done_9),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_9),
    .up_tx_rate (up_tx_rate_9),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_9),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_9),
    .up_tx_sel (up_tx_sel_9),
    .up_tx_enb (up_tx_enb_9),
    .up_tx_addr (up_tx_addr_9),
    .up_tx_wr (up_tx_wr_9),
    .up_tx_wdata (up_tx_wdata_9),
    .up_tx_rdata (up_tx_rdata_9),
    .up_tx_ready (up_tx_ready_9));
  end else begin
  assign rx_out_clk_9 = 1'd0;
  assign rx_charisk_9 = 4'd0;
  assign rx_disperr_9 = 4'd0;
  assign rx_notintable_9 = 4'd0;
  assign rx_data_9 = 32'd0;
  assign tx_9_p = 1'd0;
  assign tx_9_n = 1'd0;
  assign tx_out_clk_9 = 1'd0;
  assign up_es_rdata_9 = 16'd0;
  assign up_es_ready_9 = 1'd0;
  assign up_rx_pll_locked_9 = 1'd0;
  assign up_rx_rst_done_9 = 1'd0;
  assign up_rx_rdata_9 = 16'd0;
  assign up_rx_ready_9 = 1'd0;
  assign up_tx_pll_locked_9 = 1'd0;
  assign up_tx_rst_done_9 = 1'd0;
  assign up_tx_rdata_9 = 16'd0;
  assign up_tx_ready_9 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 11) begin
  util_adxcvr_xch #(
    .XCVR_ID (10),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_10 (
    .qpll2ch_clk (qpll2ch_clk_8),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_8),
    .qpll2ch_locked (qpll2ch_locked_8),
    .cpll_ref_clk (cpll_ref_clk_10),
    .up_cpll_rst (up_cpll_rst_10),
    .rx_p (rx_10_p),
    .rx_n (rx_10_n),
    .rx_out_clk (rx_out_clk_10),
    .rx_clk (rx_clk_10),
    .rx_charisk (rx_charisk_10),
    .rx_disperr (rx_disperr_10),
    .rx_notintable (rx_notintable_10),
    .rx_data (rx_data_10),
    .rx_calign (rx_calign_10),
    .tx_p (tx_10_p),
    .tx_n (tx_10_n),
    .tx_out_clk (tx_out_clk_10),
    .tx_clk (tx_clk_10),
    .tx_charisk (tx_charisk_10),
    .tx_data (tx_data_10),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_10),
    .up_es_enb (up_es_enb_10),
    .up_es_addr (up_es_addr_10),
    .up_es_wr (up_es_wr_10),
    .up_es_wdata (up_es_wdata_10),
    .up_es_rdata (up_es_rdata_10),
    .up_es_ready (up_es_ready_10),
    .up_rx_pll_locked (up_rx_pll_locked_10),
    .up_rx_rst (up_rx_rst_10),
    .up_rx_user_ready (up_rx_user_ready_10),
    .up_rx_rst_done (up_rx_rst_done_10),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_10),
    .up_rx_rate (up_rx_rate_10),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_10),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_10),
    .up_rx_sel (up_rx_sel_10),
    .up_rx_enb (up_rx_enb_10),
    .up_rx_addr (up_rx_addr_10),
    .up_rx_wr (up_rx_wr_10),
    .up_rx_wdata (up_rx_wdata_10),
    .up_rx_rdata (up_rx_rdata_10),
    .up_rx_ready (up_rx_ready_10),
    .up_tx_pll_locked (up_tx_pll_locked_10),
    .up_tx_rst (up_tx_rst_10),
    .up_tx_user_ready (up_tx_user_ready_10),
    .up_tx_rst_done (up_tx_rst_done_10),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_10),
    .up_tx_rate (up_tx_rate_10),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_10),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_10),
    .up_tx_sel (up_tx_sel_10),
    .up_tx_enb (up_tx_enb_10),
    .up_tx_addr (up_tx_addr_10),
    .up_tx_wr (up_tx_wr_10),
    .up_tx_wdata (up_tx_wdata_10),
    .up_tx_rdata (up_tx_rdata_10),
    .up_tx_ready (up_tx_ready_10));
  end else begin
  assign rx_out_clk_10 = 1'd0;
  assign rx_charisk_10 = 4'd0;
  assign rx_disperr_10 = 4'd0;
  assign rx_notintable_10 = 4'd0;
  assign rx_data_10 = 32'd0;
  assign tx_10_p = 1'd0;
  assign tx_10_n = 1'd0;
  assign tx_out_clk_10 = 1'd0;
  assign up_es_rdata_10 = 16'd0;
  assign up_es_ready_10 = 1'd0;
  assign up_rx_pll_locked_10 = 1'd0;
  assign up_rx_rst_done_10 = 1'd0;
  assign up_rx_rdata_10 = 16'd0;
  assign up_rx_ready_10 = 1'd0;
  assign up_tx_pll_locked_10 = 1'd0;
  assign up_tx_rst_done_10 = 1'd0;
  assign up_tx_rdata_10 = 16'd0;
  assign up_tx_ready_10 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 12) begin
  util_adxcvr_xch #(
    .XCVR_ID (11),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_11 (
    .qpll2ch_clk (qpll2ch_clk_8),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_8),
    .qpll2ch_locked (qpll2ch_locked_8),
    .cpll_ref_clk (cpll_ref_clk_11),
    .up_cpll_rst (up_cpll_rst_11),
    .rx_p (rx_11_p),
    .rx_n (rx_11_n),
    .rx_out_clk (rx_out_clk_11),
    .rx_clk (rx_clk_11),
    .rx_charisk (rx_charisk_11),
    .rx_disperr (rx_disperr_11),
    .rx_notintable (rx_notintable_11),
    .rx_data (rx_data_11),
    .rx_calign (rx_calign_11),
    .tx_p (tx_11_p),
    .tx_n (tx_11_n),
    .tx_out_clk (tx_out_clk_11),
    .tx_clk (tx_clk_11),
    .tx_charisk (tx_charisk_11),
    .tx_data (tx_data_11),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_11),
    .up_es_enb (up_es_enb_11),
    .up_es_addr (up_es_addr_11),
    .up_es_wr (up_es_wr_11),
    .up_es_wdata (up_es_wdata_11),
    .up_es_rdata (up_es_rdata_11),
    .up_es_ready (up_es_ready_11),
    .up_rx_pll_locked (up_rx_pll_locked_11),
    .up_rx_rst (up_rx_rst_11),
    .up_rx_user_ready (up_rx_user_ready_11),
    .up_rx_rst_done (up_rx_rst_done_11),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_11),
    .up_rx_rate (up_rx_rate_11),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_11),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_11),
    .up_rx_sel (up_rx_sel_11),
    .up_rx_enb (up_rx_enb_11),
    .up_rx_addr (up_rx_addr_11),
    .up_rx_wr (up_rx_wr_11),
    .up_rx_wdata (up_rx_wdata_11),
    .up_rx_rdata (up_rx_rdata_11),
    .up_rx_ready (up_rx_ready_11),
    .up_tx_pll_locked (up_tx_pll_locked_11),
    .up_tx_rst (up_tx_rst_11),
    .up_tx_user_ready (up_tx_user_ready_11),
    .up_tx_rst_done (up_tx_rst_done_11),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_11),
    .up_tx_rate (up_tx_rate_11),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_11),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_11),
    .up_tx_sel (up_tx_sel_11),
    .up_tx_enb (up_tx_enb_11),
    .up_tx_addr (up_tx_addr_11),
    .up_tx_wr (up_tx_wr_11),
    .up_tx_wdata (up_tx_wdata_11),
    .up_tx_rdata (up_tx_rdata_11),
    .up_tx_ready (up_tx_ready_11));
  end else begin
  assign rx_out_clk_11 = 1'd0;
  assign rx_charisk_11 = 4'd0;
  assign rx_disperr_11 = 4'd0;
  assign rx_notintable_11 = 4'd0;
  assign rx_data_11 = 32'd0;
  assign tx_11_p = 1'd0;
  assign tx_11_n = 1'd0;
  assign tx_out_clk_11 = 1'd0;
  assign up_es_rdata_11 = 16'd0;
  assign up_es_ready_11 = 1'd0;
  assign up_rx_pll_locked_11 = 1'd0;
  assign up_rx_rst_done_11 = 1'd0;
  assign up_rx_rdata_11 = 16'd0;
  assign up_rx_ready_11 = 1'd0;
  assign up_tx_pll_locked_11 = 1'd0;
  assign up_tx_rst_done_11 = 1'd0;
  assign up_tx_rdata_11 = 16'd0;
  assign up_tx_ready_11 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 13) begin
  util_adxcvr_xcm #(
    .XCVR_ID (12),
    .XCVR_TYPE (XCVR_TYPE),
    .QPLL_REFCLK_DIV (QPLL_REFCLK_DIV),
    .QPLL_FBDIV_RATIO (QPLL_FBDIV_RATIO),
    .QPLL_CFG (QPLL_CFG),
    .QPLL_FBDIV (QPLL_FBDIV))
  i_xcm_12 (
    .qpll_ref_clk (qpll_ref_clk_12),
    .qpll2ch_clk (qpll2ch_clk_12),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_12),
    .qpll2ch_locked (qpll2ch_locked_12),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_qpll_rst (up_qpll_rst_12),
    .up_cm_sel (up_cm_sel_12),
    .up_cm_enb (up_cm_enb_12),
    .up_cm_addr (up_cm_addr_12),
    .up_cm_wr (up_cm_wr_12),
    .up_cm_wdata (up_cm_wdata_12),
    .up_cm_rdata (up_cm_rdata_12),
    .up_cm_ready (up_cm_ready_12));
  end else begin
  assign qpll2ch_clk_12 = 1'd0;
  assign qpll2ch_ref_clk_12 = 1'd0;
  assign qpll2ch_locked_12 = 1'd0;
  assign up_cm_rdata_12 = 16'd0;
  assign up_cm_ready_12 = 1'd0;
  end
  endgenerate

  generate
  if (NUM_OF_LANES >= 13) begin
  util_adxcvr_xch #(
    .XCVR_ID (12),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_12 (
    .qpll2ch_clk (qpll2ch_clk_12),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_12),
    .qpll2ch_locked (qpll2ch_locked_12),
    .cpll_ref_clk (cpll_ref_clk_12),
    .up_cpll_rst (up_cpll_rst_12),
    .rx_p (rx_12_p),
    .rx_n (rx_12_n),
    .rx_out_clk (rx_out_clk_12),
    .rx_clk (rx_clk_12),
    .rx_charisk (rx_charisk_12),
    .rx_disperr (rx_disperr_12),
    .rx_notintable (rx_notintable_12),
    .rx_data (rx_data_12),
    .rx_calign (rx_calign_12),
    .tx_p (tx_12_p),
    .tx_n (tx_12_n),
    .tx_out_clk (tx_out_clk_12),
    .tx_clk (tx_clk_12),
    .tx_charisk (tx_charisk_12),
    .tx_data (tx_data_12),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_12),
    .up_es_enb (up_es_enb_12),
    .up_es_addr (up_es_addr_12),
    .up_es_wr (up_es_wr_12),
    .up_es_wdata (up_es_wdata_12),
    .up_es_rdata (up_es_rdata_12),
    .up_es_ready (up_es_ready_12),
    .up_rx_pll_locked (up_rx_pll_locked_12),
    .up_rx_rst (up_rx_rst_12),
    .up_rx_user_ready (up_rx_user_ready_12),
    .up_rx_rst_done (up_rx_rst_done_12),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_12),
    .up_rx_rate (up_rx_rate_12),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_12),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_12),
    .up_rx_sel (up_rx_sel_12),
    .up_rx_enb (up_rx_enb_12),
    .up_rx_addr (up_rx_addr_12),
    .up_rx_wr (up_rx_wr_12),
    .up_rx_wdata (up_rx_wdata_12),
    .up_rx_rdata (up_rx_rdata_12),
    .up_rx_ready (up_rx_ready_12),
    .up_tx_pll_locked (up_tx_pll_locked_12),
    .up_tx_rst (up_tx_rst_12),
    .up_tx_user_ready (up_tx_user_ready_12),
    .up_tx_rst_done (up_tx_rst_done_12),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_12),
    .up_tx_rate (up_tx_rate_12),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_12),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_12),
    .up_tx_sel (up_tx_sel_12),
    .up_tx_enb (up_tx_enb_12),
    .up_tx_addr (up_tx_addr_12),
    .up_tx_wr (up_tx_wr_12),
    .up_tx_wdata (up_tx_wdata_12),
    .up_tx_rdata (up_tx_rdata_12),
    .up_tx_ready (up_tx_ready_12));
  end else begin
  assign rx_out_clk_12 = 1'd0;
  assign rx_charisk_12 = 4'd0;
  assign rx_disperr_12 = 4'd0;
  assign rx_notintable_12 = 4'd0;
  assign rx_data_12 = 32'd0;
  assign tx_12_p = 1'd0;
  assign tx_12_n = 1'd0;
  assign tx_out_clk_12 = 1'd0;
  assign up_es_rdata_12 = 16'd0;
  assign up_es_ready_12 = 1'd0;
  assign up_rx_pll_locked_12 = 1'd0;
  assign up_rx_rst_done_12 = 1'd0;
  assign up_rx_rdata_12 = 16'd0;
  assign up_rx_ready_12 = 1'd0;
  assign up_tx_pll_locked_12 = 1'd0;
  assign up_tx_rst_done_12 = 1'd0;
  assign up_tx_rdata_12 = 16'd0;
  assign up_tx_ready_12 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 14) begin
  util_adxcvr_xch #(
    .XCVR_ID (13),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_13 (
    .qpll2ch_clk (qpll2ch_clk_12),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_12),
    .qpll2ch_locked (qpll2ch_locked_12),
    .cpll_ref_clk (cpll_ref_clk_13),
    .up_cpll_rst (up_cpll_rst_13),
    .rx_p (rx_13_p),
    .rx_n (rx_13_n),
    .rx_out_clk (rx_out_clk_13),
    .rx_clk (rx_clk_13),
    .rx_charisk (rx_charisk_13),
    .rx_disperr (rx_disperr_13),
    .rx_notintable (rx_notintable_13),
    .rx_data (rx_data_13),
    .rx_calign (rx_calign_13),
    .tx_p (tx_13_p),
    .tx_n (tx_13_n),
    .tx_out_clk (tx_out_clk_13),
    .tx_clk (tx_clk_13),
    .tx_charisk (tx_charisk_13),
    .tx_data (tx_data_13),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_13),
    .up_es_enb (up_es_enb_13),
    .up_es_addr (up_es_addr_13),
    .up_es_wr (up_es_wr_13),
    .up_es_wdata (up_es_wdata_13),
    .up_es_rdata (up_es_rdata_13),
    .up_es_ready (up_es_ready_13),
    .up_rx_pll_locked (up_rx_pll_locked_13),
    .up_rx_rst (up_rx_rst_13),
    .up_rx_user_ready (up_rx_user_ready_13),
    .up_rx_rst_done (up_rx_rst_done_13),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_13),
    .up_rx_rate (up_rx_rate_13),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_13),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_13),
    .up_rx_sel (up_rx_sel_13),
    .up_rx_enb (up_rx_enb_13),
    .up_rx_addr (up_rx_addr_13),
    .up_rx_wr (up_rx_wr_13),
    .up_rx_wdata (up_rx_wdata_13),
    .up_rx_rdata (up_rx_rdata_13),
    .up_rx_ready (up_rx_ready_13),
    .up_tx_pll_locked (up_tx_pll_locked_13),
    .up_tx_rst (up_tx_rst_13),
    .up_tx_user_ready (up_tx_user_ready_13),
    .up_tx_rst_done (up_tx_rst_done_13),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_13),
    .up_tx_rate (up_tx_rate_13),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_13),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_13),
    .up_tx_sel (up_tx_sel_13),
    .up_tx_enb (up_tx_enb_13),
    .up_tx_addr (up_tx_addr_13),
    .up_tx_wr (up_tx_wr_13),
    .up_tx_wdata (up_tx_wdata_13),
    .up_tx_rdata (up_tx_rdata_13),
    .up_tx_ready (up_tx_ready_13));
  end else begin
  assign rx_out_clk_13 = 1'd0;
  assign rx_charisk_13 = 4'd0;
  assign rx_disperr_13 = 4'd0;
  assign rx_notintable_13 = 4'd0;
  assign rx_data_13 = 32'd0;
  assign tx_13_p = 1'd0;
  assign tx_13_n = 1'd0;
  assign tx_out_clk_13 = 1'd0;
  assign up_es_rdata_13 = 16'd0;
  assign up_es_ready_13 = 1'd0;
  assign up_rx_pll_locked_13 = 1'd0;
  assign up_rx_rst_done_13 = 1'd0;
  assign up_rx_rdata_13 = 16'd0;
  assign up_rx_ready_13 = 1'd0;
  assign up_tx_pll_locked_13 = 1'd0;
  assign up_tx_rst_done_13 = 1'd0;
  assign up_tx_rdata_13 = 16'd0;
  assign up_tx_ready_13 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 15) begin
  util_adxcvr_xch #(
    .XCVR_ID (14),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_14 (
    .qpll2ch_clk (qpll2ch_clk_12),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_12),
    .qpll2ch_locked (qpll2ch_locked_12),
    .cpll_ref_clk (cpll_ref_clk_14),
    .up_cpll_rst (up_cpll_rst_14),
    .rx_p (rx_14_p),
    .rx_n (rx_14_n),
    .rx_out_clk (rx_out_clk_14),
    .rx_clk (rx_clk_14),
    .rx_charisk (rx_charisk_14),
    .rx_disperr (rx_disperr_14),
    .rx_notintable (rx_notintable_14),
    .rx_data (rx_data_14),
    .rx_calign (rx_calign_14),
    .tx_p (tx_14_p),
    .tx_n (tx_14_n),
    .tx_out_clk (tx_out_clk_14),
    .tx_clk (tx_clk_14),
    .tx_charisk (tx_charisk_14),
    .tx_data (tx_data_14),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_14),
    .up_es_enb (up_es_enb_14),
    .up_es_addr (up_es_addr_14),
    .up_es_wr (up_es_wr_14),
    .up_es_wdata (up_es_wdata_14),
    .up_es_rdata (up_es_rdata_14),
    .up_es_ready (up_es_ready_14),
    .up_rx_pll_locked (up_rx_pll_locked_14),
    .up_rx_rst (up_rx_rst_14),
    .up_rx_user_ready (up_rx_user_ready_14),
    .up_rx_rst_done (up_rx_rst_done_14),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_14),
    .up_rx_rate (up_rx_rate_14),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_14),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_14),
    .up_rx_sel (up_rx_sel_14),
    .up_rx_enb (up_rx_enb_14),
    .up_rx_addr (up_rx_addr_14),
    .up_rx_wr (up_rx_wr_14),
    .up_rx_wdata (up_rx_wdata_14),
    .up_rx_rdata (up_rx_rdata_14),
    .up_rx_ready (up_rx_ready_14),
    .up_tx_pll_locked (up_tx_pll_locked_14),
    .up_tx_rst (up_tx_rst_14),
    .up_tx_user_ready (up_tx_user_ready_14),
    .up_tx_rst_done (up_tx_rst_done_14),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_14),
    .up_tx_rate (up_tx_rate_14),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_14),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_14),
    .up_tx_sel (up_tx_sel_14),
    .up_tx_enb (up_tx_enb_14),
    .up_tx_addr (up_tx_addr_14),
    .up_tx_wr (up_tx_wr_14),
    .up_tx_wdata (up_tx_wdata_14),
    .up_tx_rdata (up_tx_rdata_14),
    .up_tx_ready (up_tx_ready_14));
  end else begin
  assign rx_out_clk_14 = 1'd0;
  assign rx_charisk_14 = 4'd0;
  assign rx_disperr_14 = 4'd0;
  assign rx_notintable_14 = 4'd0;
  assign rx_data_14 = 32'd0;
  assign tx_14_p = 1'd0;
  assign tx_14_n = 1'd0;
  assign tx_out_clk_14 = 1'd0;
  assign up_es_rdata_14 = 16'd0;
  assign up_es_ready_14 = 1'd0;
  assign up_rx_pll_locked_14 = 1'd0;
  assign up_rx_rst_done_14 = 1'd0;
  assign up_rx_rdata_14 = 16'd0;
  assign up_rx_ready_14 = 1'd0;
  assign up_tx_pll_locked_14 = 1'd0;
  assign up_tx_rst_done_14 = 1'd0;
  assign up_tx_rdata_14 = 16'd0;
  assign up_tx_ready_14 = 1'd0;
  end
  endgenerate


  generate
  if (NUM_OF_LANES >= 16) begin
  util_adxcvr_xch #(
    .XCVR_ID (15),
    .XCVR_TYPE (XCVR_TYPE),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_4_5 (CPLL_FBDIV_4_5),
    .TX_OUT_DIV (TX_OUT_DIV),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .RX_OUT_DIV (RX_OUT_DIV),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_PMA_CFG (RX_PMA_CFG),
    .RX_CDR_CFG (RX_CDR_CFG))
  i_xch_15 (
    .qpll2ch_clk (qpll2ch_clk_12),
    .qpll2ch_ref_clk (qpll2ch_ref_clk_12),
    .qpll2ch_locked (qpll2ch_locked_12),
    .cpll_ref_clk (cpll_ref_clk_15),
    .up_cpll_rst (up_cpll_rst_15),
    .rx_p (rx_15_p),
    .rx_n (rx_15_n),
    .rx_out_clk (rx_out_clk_15),
    .rx_clk (rx_clk_15),
    .rx_charisk (rx_charisk_15),
    .rx_disperr (rx_disperr_15),
    .rx_notintable (rx_notintable_15),
    .rx_data (rx_data_15),
    .rx_calign (rx_calign_15),
    .tx_p (tx_15_p),
    .tx_n (tx_15_n),
    .tx_out_clk (tx_out_clk_15),
    .tx_clk (tx_clk_15),
    .tx_charisk (tx_charisk_15),
    .tx_data (tx_data_15),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_sel (up_es_sel_15),
    .up_es_enb (up_es_enb_15),
    .up_es_addr (up_es_addr_15),
    .up_es_wr (up_es_wr_15),
    .up_es_wdata (up_es_wdata_15),
    .up_es_rdata (up_es_rdata_15),
    .up_es_ready (up_es_ready_15),
    .up_rx_pll_locked (up_rx_pll_locked_15),
    .up_rx_rst (up_rx_rst_15),
    .up_rx_user_ready (up_rx_user_ready_15),
    .up_rx_rst_done (up_rx_rst_done_15),
    .up_rx_lpm_dfe_n (up_rx_lpm_dfe_n_15),
    .up_rx_rate (up_rx_rate_15),
    .up_rx_sys_clk_sel (up_rx_sys_clk_sel_15),
    .up_rx_out_clk_sel (up_rx_out_clk_sel_15),
    .up_rx_sel (up_rx_sel_15),
    .up_rx_enb (up_rx_enb_15),
    .up_rx_addr (up_rx_addr_15),
    .up_rx_wr (up_rx_wr_15),
    .up_rx_wdata (up_rx_wdata_15),
    .up_rx_rdata (up_rx_rdata_15),
    .up_rx_ready (up_rx_ready_15),
    .up_tx_pll_locked (up_tx_pll_locked_15),
    .up_tx_rst (up_tx_rst_15),
    .up_tx_user_ready (up_tx_user_ready_15),
    .up_tx_rst_done (up_tx_rst_done_15),
    .up_tx_lpm_dfe_n (up_tx_lpm_dfe_n_15),
    .up_tx_rate (up_tx_rate_15),
    .up_tx_sys_clk_sel (up_tx_sys_clk_sel_15),
    .up_tx_out_clk_sel (up_tx_out_clk_sel_15),
    .up_tx_sel (up_tx_sel_15),
    .up_tx_enb (up_tx_enb_15),
    .up_tx_addr (up_tx_addr_15),
    .up_tx_wr (up_tx_wr_15),
    .up_tx_wdata (up_tx_wdata_15),
    .up_tx_rdata (up_tx_rdata_15),
    .up_tx_ready (up_tx_ready_15));
  end else begin
  assign rx_out_clk_15 = 1'd0;
  assign rx_charisk_15 = 4'd0;
  assign rx_disperr_15 = 4'd0;
  assign rx_notintable_15 = 4'd0;
  assign rx_data_15 = 32'd0;
  assign tx_15_p = 1'd0;
  assign tx_15_n = 1'd0;
  assign tx_out_clk_15 = 1'd0;
  assign up_es_rdata_15 = 16'd0;
  assign up_es_ready_15 = 1'd0;
  assign up_rx_pll_locked_15 = 1'd0;
  assign up_rx_rst_done_15 = 1'd0;
  assign up_rx_rdata_15 = 16'd0;
  assign up_rx_ready_15 = 1'd0;
  assign up_tx_pll_locked_15 = 1'd0;
  assign up_tx_rst_done_15 = 1'd0;
  assign up_tx_rdata_15 = 16'd0;
  assign up_tx_ready_15 = 1'd0;
  end
  endgenerate

endmodule

// ***************************************************************************
// ***************************************************************************


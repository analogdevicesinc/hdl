// ***************************************************************************
// ***************************************************************************
// Copyright 2014 - 2017 (c) Analog Devices, Inc. All rights reserved.
//
// Each core or library found in this collection may have its own licensing terms. 
// The user should keep this in in mind while exploring these cores. 
//
// Redistribution and use in source and binary forms,
// with or without modification of this file, are permitted under the terms of either
//  (at the option of the user):
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory, or at:
// https://www.gnu.org/licenses/old-licenses/gpl-2.0.en.html
//
// OR
//
//   2.  An ADI specific BSD license as noted in the top level directory, or on-line at:
// https://github.com/analogdevicesinc/hdl/blob/dev/LICENSE
//
// ***************************************************************************
// ***************************************************************************
// AUTO GENERATED BY axi_adxcvr.pl, DO NOT MODIFY!

`timescale 1ns/1ps

module axi_adxcvr #(

  // parameters

  parameter   integer ID = 0,
  parameter   integer NUM_OF_LANES = 8,
  parameter   integer GTH_OR_GTX_N = 0,
  parameter   integer TX_OR_RX_N = 0,
  parameter   integer QPLL_ENABLE = 1,
  parameter           LPM_OR_DFE_N = 1,
  parameter   [ 2:0]  RATE = 3'd0,
  parameter   [ 1:0]  SYS_CLK_SEL = 2'd3,
  parameter   [ 2:0]  OUT_CLK_SEL = 3'd4) (

  output  [ 7:0]  up_cm_sel_0,
  output          up_cm_enb_0,
  output  [11:0]  up_cm_addr_0,
  output          up_cm_wr_0,
  output  [15:0]  up_cm_wdata_0,
  input   [15:0]  up_cm_rdata_0,
  input           up_cm_ready_0,

  output  [ 7:0]  up_es_sel_0,
  output          up_es_enb_0,
  output  [11:0]  up_es_addr_0,
  output          up_es_wr_0,
  output  [15:0]  up_es_wdata_0,
  input   [15:0]  up_es_rdata_0,
  input           up_es_ready_0,

  input           up_ch_pll_locked_0,
  output          up_ch_rst_0,
  output          up_ch_user_ready_0,
  input           up_ch_rst_done_0,
  output          up_ch_lpm_dfe_n_0,
  output  [ 2:0]  up_ch_rate_0,
  output  [ 1:0]  up_ch_sys_clk_sel_0,
  output  [ 2:0]  up_ch_out_clk_sel_0,
  output  [ 7:0]  up_ch_sel_0,
  output          up_ch_enb_0,
  output  [11:0]  up_ch_addr_0,
  output          up_ch_wr_0,
  output  [15:0]  up_ch_wdata_0,
  input   [15:0]  up_ch_rdata_0,
  input           up_ch_ready_0,

  output  [ 7:0]  up_es_sel_1,
  output          up_es_enb_1,
  output  [11:0]  up_es_addr_1,
  output          up_es_wr_1,
  output  [15:0]  up_es_wdata_1,
  input   [15:0]  up_es_rdata_1,
  input           up_es_ready_1,

  input           up_ch_pll_locked_1,
  output          up_ch_rst_1,
  output          up_ch_user_ready_1,
  input           up_ch_rst_done_1,
  output          up_ch_lpm_dfe_n_1,
  output  [ 2:0]  up_ch_rate_1,
  output  [ 1:0]  up_ch_sys_clk_sel_1,
  output  [ 2:0]  up_ch_out_clk_sel_1,
  output  [ 7:0]  up_ch_sel_1,
  output          up_ch_enb_1,
  output  [11:0]  up_ch_addr_1,
  output          up_ch_wr_1,
  output  [15:0]  up_ch_wdata_1,
  input   [15:0]  up_ch_rdata_1,
  input           up_ch_ready_1,

  output  [ 7:0]  up_es_sel_2,
  output          up_es_enb_2,
  output  [11:0]  up_es_addr_2,
  output          up_es_wr_2,
  output  [15:0]  up_es_wdata_2,
  input   [15:0]  up_es_rdata_2,
  input           up_es_ready_2,

  input           up_ch_pll_locked_2,
  output          up_ch_rst_2,
  output          up_ch_user_ready_2,
  input           up_ch_rst_done_2,
  output          up_ch_lpm_dfe_n_2,
  output  [ 2:0]  up_ch_rate_2,
  output  [ 1:0]  up_ch_sys_clk_sel_2,
  output  [ 2:0]  up_ch_out_clk_sel_2,
  output  [ 7:0]  up_ch_sel_2,
  output          up_ch_enb_2,
  output  [11:0]  up_ch_addr_2,
  output          up_ch_wr_2,
  output  [15:0]  up_ch_wdata_2,
  input   [15:0]  up_ch_rdata_2,
  input           up_ch_ready_2,

  output  [ 7:0]  up_es_sel_3,
  output          up_es_enb_3,
  output  [11:0]  up_es_addr_3,
  output          up_es_wr_3,
  output  [15:0]  up_es_wdata_3,
  input   [15:0]  up_es_rdata_3,
  input           up_es_ready_3,

  input           up_ch_pll_locked_3,
  output          up_ch_rst_3,
  output          up_ch_user_ready_3,
  input           up_ch_rst_done_3,
  output          up_ch_lpm_dfe_n_3,
  output  [ 2:0]  up_ch_rate_3,
  output  [ 1:0]  up_ch_sys_clk_sel_3,
  output  [ 2:0]  up_ch_out_clk_sel_3,
  output  [ 7:0]  up_ch_sel_3,
  output          up_ch_enb_3,
  output  [11:0]  up_ch_addr_3,
  output          up_ch_wr_3,
  output  [15:0]  up_ch_wdata_3,
  input   [15:0]  up_ch_rdata_3,
  input           up_ch_ready_3,

  output  [ 7:0]  up_cm_sel_4,
  output          up_cm_enb_4,
  output  [11:0]  up_cm_addr_4,
  output          up_cm_wr_4,
  output  [15:0]  up_cm_wdata_4,
  input   [15:0]  up_cm_rdata_4,
  input           up_cm_ready_4,

  output  [ 7:0]  up_es_sel_4,
  output          up_es_enb_4,
  output  [11:0]  up_es_addr_4,
  output          up_es_wr_4,
  output  [15:0]  up_es_wdata_4,
  input   [15:0]  up_es_rdata_4,
  input           up_es_ready_4,

  input           up_ch_pll_locked_4,
  output          up_ch_rst_4,
  output          up_ch_user_ready_4,
  input           up_ch_rst_done_4,
  output          up_ch_lpm_dfe_n_4,
  output  [ 2:0]  up_ch_rate_4,
  output  [ 1:0]  up_ch_sys_clk_sel_4,
  output  [ 2:0]  up_ch_out_clk_sel_4,
  output  [ 7:0]  up_ch_sel_4,
  output          up_ch_enb_4,
  output  [11:0]  up_ch_addr_4,
  output          up_ch_wr_4,
  output  [15:0]  up_ch_wdata_4,
  input   [15:0]  up_ch_rdata_4,
  input           up_ch_ready_4,

  output  [ 7:0]  up_es_sel_5,
  output          up_es_enb_5,
  output  [11:0]  up_es_addr_5,
  output          up_es_wr_5,
  output  [15:0]  up_es_wdata_5,
  input   [15:0]  up_es_rdata_5,
  input           up_es_ready_5,

  input           up_ch_pll_locked_5,
  output          up_ch_rst_5,
  output          up_ch_user_ready_5,
  input           up_ch_rst_done_5,
  output          up_ch_lpm_dfe_n_5,
  output  [ 2:0]  up_ch_rate_5,
  output  [ 1:0]  up_ch_sys_clk_sel_5,
  output  [ 2:0]  up_ch_out_clk_sel_5,
  output  [ 7:0]  up_ch_sel_5,
  output          up_ch_enb_5,
  output  [11:0]  up_ch_addr_5,
  output          up_ch_wr_5,
  output  [15:0]  up_ch_wdata_5,
  input   [15:0]  up_ch_rdata_5,
  input           up_ch_ready_5,

  output  [ 7:0]  up_es_sel_6,
  output          up_es_enb_6,
  output  [11:0]  up_es_addr_6,
  output          up_es_wr_6,
  output  [15:0]  up_es_wdata_6,
  input   [15:0]  up_es_rdata_6,
  input           up_es_ready_6,

  input           up_ch_pll_locked_6,
  output          up_ch_rst_6,
  output          up_ch_user_ready_6,
  input           up_ch_rst_done_6,
  output          up_ch_lpm_dfe_n_6,
  output  [ 2:0]  up_ch_rate_6,
  output  [ 1:0]  up_ch_sys_clk_sel_6,
  output  [ 2:0]  up_ch_out_clk_sel_6,
  output  [ 7:0]  up_ch_sel_6,
  output          up_ch_enb_6,
  output  [11:0]  up_ch_addr_6,
  output          up_ch_wr_6,
  output  [15:0]  up_ch_wdata_6,
  input   [15:0]  up_ch_rdata_6,
  input           up_ch_ready_6,

  output  [ 7:0]  up_es_sel_7,
  output          up_es_enb_7,
  output  [11:0]  up_es_addr_7,
  output          up_es_wr_7,
  output  [15:0]  up_es_wdata_7,
  input   [15:0]  up_es_rdata_7,
  input           up_es_ready_7,

  input           up_ch_pll_locked_7,
  output          up_ch_rst_7,
  output          up_ch_user_ready_7,
  input           up_ch_rst_done_7,
  output          up_ch_lpm_dfe_n_7,
  output  [ 2:0]  up_ch_rate_7,
  output  [ 1:0]  up_ch_sys_clk_sel_7,
  output  [ 2:0]  up_ch_out_clk_sel_7,
  output  [ 7:0]  up_ch_sel_7,
  output          up_ch_enb_7,
  output  [11:0]  up_ch_addr_7,
  output          up_ch_wr_7,
  output  [15:0]  up_ch_wdata_7,
  input   [15:0]  up_ch_rdata_7,
  input           up_ch_ready_7,

  output  [ 7:0]  up_cm_sel_8,
  output          up_cm_enb_8,
  output  [11:0]  up_cm_addr_8,
  output          up_cm_wr_8,
  output  [15:0]  up_cm_wdata_8,
  input   [15:0]  up_cm_rdata_8,
  input           up_cm_ready_8,

  output  [ 7:0]  up_es_sel_8,
  output          up_es_enb_8,
  output  [11:0]  up_es_addr_8,
  output          up_es_wr_8,
  output  [15:0]  up_es_wdata_8,
  input   [15:0]  up_es_rdata_8,
  input           up_es_ready_8,

  input           up_ch_pll_locked_8,
  output          up_ch_rst_8,
  output          up_ch_user_ready_8,
  input           up_ch_rst_done_8,
  output          up_ch_lpm_dfe_n_8,
  output  [ 2:0]  up_ch_rate_8,
  output  [ 1:0]  up_ch_sys_clk_sel_8,
  output  [ 2:0]  up_ch_out_clk_sel_8,
  output  [ 7:0]  up_ch_sel_8,
  output          up_ch_enb_8,
  output  [11:0]  up_ch_addr_8,
  output          up_ch_wr_8,
  output  [15:0]  up_ch_wdata_8,
  input   [15:0]  up_ch_rdata_8,
  input           up_ch_ready_8,

  output  [ 7:0]  up_es_sel_9,
  output          up_es_enb_9,
  output  [11:0]  up_es_addr_9,
  output          up_es_wr_9,
  output  [15:0]  up_es_wdata_9,
  input   [15:0]  up_es_rdata_9,
  input           up_es_ready_9,

  input           up_ch_pll_locked_9,
  output          up_ch_rst_9,
  output          up_ch_user_ready_9,
  input           up_ch_rst_done_9,
  output          up_ch_lpm_dfe_n_9,
  output  [ 2:0]  up_ch_rate_9,
  output  [ 1:0]  up_ch_sys_clk_sel_9,
  output  [ 2:0]  up_ch_out_clk_sel_9,
  output  [ 7:0]  up_ch_sel_9,
  output          up_ch_enb_9,
  output  [11:0]  up_ch_addr_9,
  output          up_ch_wr_9,
  output  [15:0]  up_ch_wdata_9,
  input   [15:0]  up_ch_rdata_9,
  input           up_ch_ready_9,

  output  [ 7:0]  up_es_sel_10,
  output          up_es_enb_10,
  output  [11:0]  up_es_addr_10,
  output          up_es_wr_10,
  output  [15:0]  up_es_wdata_10,
  input   [15:0]  up_es_rdata_10,
  input           up_es_ready_10,

  input           up_ch_pll_locked_10,
  output          up_ch_rst_10,
  output          up_ch_user_ready_10,
  input           up_ch_rst_done_10,
  output          up_ch_lpm_dfe_n_10,
  output  [ 2:0]  up_ch_rate_10,
  output  [ 1:0]  up_ch_sys_clk_sel_10,
  output  [ 2:0]  up_ch_out_clk_sel_10,
  output  [ 7:0]  up_ch_sel_10,
  output          up_ch_enb_10,
  output  [11:0]  up_ch_addr_10,
  output          up_ch_wr_10,
  output  [15:0]  up_ch_wdata_10,
  input   [15:0]  up_ch_rdata_10,
  input           up_ch_ready_10,

  output  [ 7:0]  up_es_sel_11,
  output          up_es_enb_11,
  output  [11:0]  up_es_addr_11,
  output          up_es_wr_11,
  output  [15:0]  up_es_wdata_11,
  input   [15:0]  up_es_rdata_11,
  input           up_es_ready_11,

  input           up_ch_pll_locked_11,
  output          up_ch_rst_11,
  output          up_ch_user_ready_11,
  input           up_ch_rst_done_11,
  output          up_ch_lpm_dfe_n_11,
  output  [ 2:0]  up_ch_rate_11,
  output  [ 1:0]  up_ch_sys_clk_sel_11,
  output  [ 2:0]  up_ch_out_clk_sel_11,
  output  [ 7:0]  up_ch_sel_11,
  output          up_ch_enb_11,
  output  [11:0]  up_ch_addr_11,
  output          up_ch_wr_11,
  output  [15:0]  up_ch_wdata_11,
  input   [15:0]  up_ch_rdata_11,
  input           up_ch_ready_11,

  output  [ 7:0]  up_cm_sel_12,
  output          up_cm_enb_12,
  output  [11:0]  up_cm_addr_12,
  output          up_cm_wr_12,
  output  [15:0]  up_cm_wdata_12,
  input   [15:0]  up_cm_rdata_12,
  input           up_cm_ready_12,

  output  [ 7:0]  up_es_sel_12,
  output          up_es_enb_12,
  output  [11:0]  up_es_addr_12,
  output          up_es_wr_12,
  output  [15:0]  up_es_wdata_12,
  input   [15:0]  up_es_rdata_12,
  input           up_es_ready_12,

  input           up_ch_pll_locked_12,
  output          up_ch_rst_12,
  output          up_ch_user_ready_12,
  input           up_ch_rst_done_12,
  output          up_ch_lpm_dfe_n_12,
  output  [ 2:0]  up_ch_rate_12,
  output  [ 1:0]  up_ch_sys_clk_sel_12,
  output  [ 2:0]  up_ch_out_clk_sel_12,
  output  [ 7:0]  up_ch_sel_12,
  output          up_ch_enb_12,
  output  [11:0]  up_ch_addr_12,
  output          up_ch_wr_12,
  output  [15:0]  up_ch_wdata_12,
  input   [15:0]  up_ch_rdata_12,
  input           up_ch_ready_12,

  output  [ 7:0]  up_es_sel_13,
  output          up_es_enb_13,
  output  [11:0]  up_es_addr_13,
  output          up_es_wr_13,
  output  [15:0]  up_es_wdata_13,
  input   [15:0]  up_es_rdata_13,
  input           up_es_ready_13,

  input           up_ch_pll_locked_13,
  output          up_ch_rst_13,
  output          up_ch_user_ready_13,
  input           up_ch_rst_done_13,
  output          up_ch_lpm_dfe_n_13,
  output  [ 2:0]  up_ch_rate_13,
  output  [ 1:0]  up_ch_sys_clk_sel_13,
  output  [ 2:0]  up_ch_out_clk_sel_13,
  output  [ 7:0]  up_ch_sel_13,
  output          up_ch_enb_13,
  output  [11:0]  up_ch_addr_13,
  output          up_ch_wr_13,
  output  [15:0]  up_ch_wdata_13,
  input   [15:0]  up_ch_rdata_13,
  input           up_ch_ready_13,

  output  [ 7:0]  up_es_sel_14,
  output          up_es_enb_14,
  output  [11:0]  up_es_addr_14,
  output          up_es_wr_14,
  output  [15:0]  up_es_wdata_14,
  input   [15:0]  up_es_rdata_14,
  input           up_es_ready_14,

  input           up_ch_pll_locked_14,
  output          up_ch_rst_14,
  output          up_ch_user_ready_14,
  input           up_ch_rst_done_14,
  output          up_ch_lpm_dfe_n_14,
  output  [ 2:0]  up_ch_rate_14,
  output  [ 1:0]  up_ch_sys_clk_sel_14,
  output  [ 2:0]  up_ch_out_clk_sel_14,
  output  [ 7:0]  up_ch_sel_14,
  output          up_ch_enb_14,
  output  [11:0]  up_ch_addr_14,
  output          up_ch_wr_14,
  output  [15:0]  up_ch_wdata_14,
  input   [15:0]  up_ch_rdata_14,
  input           up_ch_ready_14,

  output  [ 7:0]  up_es_sel_15,
  output          up_es_enb_15,
  output  [11:0]  up_es_addr_15,
  output          up_es_wr_15,
  output  [15:0]  up_es_wdata_15,
  input   [15:0]  up_es_rdata_15,
  input           up_es_ready_15,

  input           up_ch_pll_locked_15,
  output          up_ch_rst_15,
  output          up_ch_user_ready_15,
  input           up_ch_rst_done_15,
  output          up_ch_lpm_dfe_n_15,
  output  [ 2:0]  up_ch_rate_15,
  output  [ 1:0]  up_ch_sys_clk_sel_15,
  output  [ 2:0]  up_ch_out_clk_sel_15,
  output  [ 7:0]  up_ch_sel_15,
  output          up_ch_enb_15,
  output  [11:0]  up_ch_addr_15,
  output          up_ch_wr_15,
  output  [15:0]  up_ch_wdata_15,
  input   [15:0]  up_ch_rdata_15,
  input           up_ch_ready_15,

  input           s_axi_aclk,
  input           s_axi_aresetn,
  output          up_status,
  output          up_pll_rst,

  input           s_axi_awvalid,
  input   [31:0]  s_axi_awaddr,
  input   [ 2:0]  s_axi_awprot,
  output          s_axi_awready,
  input           s_axi_wvalid,
  input   [31:0]  s_axi_wdata,
  input   [ 3:0]  s_axi_wstrb,
  output          s_axi_wready,
  output          s_axi_bvalid,
  output  [ 1:0]  s_axi_bresp,
  input           s_axi_bready,
  input           s_axi_arvalid,
  input   [31:0]  s_axi_araddr,
  input   [ 2:0]  s_axi_arprot,
  output          s_axi_arready,
  output          s_axi_rvalid,
  output  [ 1:0]  s_axi_rresp,
  output  [31:0]  s_axi_rdata,
  input           s_axi_rready,

  output          m_axi_awvalid,
  output  [31:0]  m_axi_awaddr,
  output  [ 2:0]  m_axi_awprot,
  input           m_axi_awready,
  output          m_axi_wvalid,
  output  [31:0]  m_axi_wdata,
  output  [ 3:0]  m_axi_wstrb,
  input           m_axi_wready,
  input           m_axi_bvalid,
  input   [ 1:0]  m_axi_bresp,
  output          m_axi_bready,
  output          m_axi_arvalid,
  output  [31:0]  m_axi_araddr,
  output  [ 2:0]  m_axi_arprot,
  input           m_axi_arready,
  input           m_axi_rvalid,
  input   [31:0]  m_axi_rdata,
  input   [ 1:0]  m_axi_rresp,
  output          m_axi_rready);

  // internal signals

  wire    [ 7:0]  up_cm_sel;
  wire            up_cm_enb;
  wire    [11:0]  up_cm_addr;
  wire            up_cm_wr;
  wire    [15:0]  up_cm_wdata;
  wire    [15:0]  up_cm_rdata_0_s;
  wire            up_cm_ready_0_s;
  wire    [15:0]  up_cm_rdata_4_s;
  wire            up_cm_ready_4_s;
  wire    [15:0]  up_cm_rdata_8_s;
  wire            up_cm_ready_8_s;
  wire    [15:0]  up_cm_rdata_12_s;
  wire            up_cm_ready_12_s;
  wire    [ 7:0]  up_es_sel;
  wire            up_es_enb;
  wire    [11:0]  up_es_addr;
  wire            up_es_wr;
  wire    [15:0]  up_es_wdata;
  wire    [15:0]  up_es_rdata_0_s;
  wire            up_es_ready_0_s;
  wire    [15:0]  up_es_rdata_1_s;
  wire            up_es_ready_1_s;
  wire    [15:0]  up_es_rdata_2_s;
  wire            up_es_ready_2_s;
  wire    [15:0]  up_es_rdata_3_s;
  wire            up_es_ready_3_s;
  wire    [15:0]  up_es_rdata_4_s;
  wire            up_es_ready_4_s;
  wire    [15:0]  up_es_rdata_5_s;
  wire            up_es_ready_5_s;
  wire    [15:0]  up_es_rdata_6_s;
  wire            up_es_ready_6_s;
  wire    [15:0]  up_es_rdata_7_s;
  wire            up_es_ready_7_s;
  wire    [15:0]  up_es_rdata_8_s;
  wire            up_es_ready_8_s;
  wire    [15:0]  up_es_rdata_9_s;
  wire            up_es_ready_9_s;
  wire    [15:0]  up_es_rdata_10_s;
  wire            up_es_ready_10_s;
  wire    [15:0]  up_es_rdata_11_s;
  wire            up_es_ready_11_s;
  wire    [15:0]  up_es_rdata_12_s;
  wire            up_es_ready_12_s;
  wire    [15:0]  up_es_rdata_13_s;
  wire            up_es_ready_13_s;
  wire    [15:0]  up_es_rdata_14_s;
  wire            up_es_ready_14_s;
  wire    [15:0]  up_es_rdata_15_s;
  wire            up_es_ready_15_s;
  wire            up_ch_rst;
  wire            up_ch_user_ready;
  wire            up_ch_lpm_dfe_n;
  wire    [ 2:0]  up_ch_rate;
  wire    [ 1:0]  up_ch_sys_clk_sel;
  wire    [ 2:0]  up_ch_out_clk_sel;
  wire            up_ch_pll_locked_0_s;
  wire            up_ch_rst_done_0_s;
  wire            up_ch_pll_locked_1_s;
  wire            up_ch_rst_done_1_s;
  wire            up_ch_pll_locked_2_s;
  wire            up_ch_rst_done_2_s;
  wire            up_ch_pll_locked_3_s;
  wire            up_ch_rst_done_3_s;
  wire            up_ch_pll_locked_4_s;
  wire            up_ch_rst_done_4_s;
  wire            up_ch_pll_locked_5_s;
  wire            up_ch_rst_done_5_s;
  wire            up_ch_pll_locked_6_s;
  wire            up_ch_rst_done_6_s;
  wire            up_ch_pll_locked_7_s;
  wire            up_ch_rst_done_7_s;
  wire            up_ch_pll_locked_8_s;
  wire            up_ch_rst_done_8_s;
  wire            up_ch_pll_locked_9_s;
  wire            up_ch_rst_done_9_s;
  wire            up_ch_pll_locked_10_s;
  wire            up_ch_rst_done_10_s;
  wire            up_ch_pll_locked_11_s;
  wire            up_ch_rst_done_11_s;
  wire            up_ch_pll_locked_12_s;
  wire            up_ch_rst_done_12_s;
  wire            up_ch_pll_locked_13_s;
  wire            up_ch_rst_done_13_s;
  wire            up_ch_pll_locked_14_s;
  wire            up_ch_rst_done_14_s;
  wire            up_ch_pll_locked_15_s;
  wire            up_ch_rst_done_15_s;
  wire    [ 7:0]  up_ch_sel;
  wire            up_ch_enb;
  wire    [11:0]  up_ch_addr;
  wire            up_ch_wr;
  wire    [15:0]  up_ch_wdata;
  wire    [15:0]  up_ch_rdata_0_s;
  wire            up_ch_ready_0_s;
  wire    [15:0]  up_ch_rdata_1_s;
  wire            up_ch_ready_1_s;
  wire    [15:0]  up_ch_rdata_2_s;
  wire            up_ch_ready_2_s;
  wire    [15:0]  up_ch_rdata_3_s;
  wire            up_ch_ready_3_s;
  wire    [15:0]  up_ch_rdata_4_s;
  wire            up_ch_ready_4_s;
  wire    [15:0]  up_ch_rdata_5_s;
  wire            up_ch_ready_5_s;
  wire    [15:0]  up_ch_rdata_6_s;
  wire            up_ch_ready_6_s;
  wire    [15:0]  up_ch_rdata_7_s;
  wire            up_ch_ready_7_s;
  wire    [15:0]  up_ch_rdata_8_s;
  wire            up_ch_ready_8_s;
  wire    [15:0]  up_ch_rdata_9_s;
  wire            up_ch_ready_9_s;
  wire    [15:0]  up_ch_rdata_10_s;
  wire            up_ch_ready_10_s;
  wire    [15:0]  up_ch_rdata_11_s;
  wire            up_ch_ready_11_s;
  wire    [15:0]  up_ch_rdata_12_s;
  wire            up_ch_ready_12_s;
  wire    [15:0]  up_ch_rdata_13_s;
  wire            up_ch_ready_13_s;
  wire    [15:0]  up_ch_rdata_14_s;
  wire            up_ch_ready_14_s;
  wire    [15:0]  up_ch_rdata_15_s;
  wire            up_ch_ready_15_s;
  wire            up_es_req;
  wire            up_es_ack;
  wire    [ 4:0]  up_es_pscale;
  wire    [ 1:0]  up_es_vrange;
  wire    [ 7:0]  up_es_vstep;
  wire    [ 7:0]  up_es_vmax;
  wire    [ 7:0]  up_es_vmin;
  wire    [11:0]  up_es_hmax;
  wire    [11:0]  up_es_hmin;
  wire    [11:0]  up_es_hstep;
  wire    [31:0]  up_es_saddr;
  wire            up_es_status;
  wire            up_rstn;
  wire            up_clk;
  wire            up_wreq;
  wire    [ 9:0]  up_waddr;
  wire    [31:0]  up_wdata;
  wire            up_wack;
  wire            up_rreq;
  wire    [ 9:0]  up_raddr;
  wire    [31:0]  up_rdata;
  wire            up_rack;

  // channel broadcast

  assign up_rstn = s_axi_aresetn;
  assign up_clk = s_axi_aclk;

  assign up_cm_sel_0 = up_cm_sel;
  assign up_cm_enb_0 = up_cm_enb;
  assign up_cm_addr_0 = up_cm_addr;
  assign up_cm_wr_0 = up_cm_wr;
  assign up_cm_wdata_0 = up_cm_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (0),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_cm_0 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_cm_sel),
    .up_enb (up_cm_enb),
    .up_rdata_in (16'd0),
    .up_ready_in (1'd1),
    .up_rdata (up_cm_rdata_0),
    .up_ready (up_cm_ready_0),
    .up_rdata_out (up_cm_rdata_0_s),
    .up_ready_out (up_cm_ready_0_s));

  assign up_es_sel_0 = up_es_sel;
  assign up_es_enb_0 = up_es_enb;
  assign up_es_addr_0 = up_es_addr;
  assign up_es_wr_0 = up_es_wr;
  assign up_es_wdata_0 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (0),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_0 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (16'd0),
    .up_ready_in (1'd1),
    .up_rdata (up_es_rdata_0),
    .up_ready (up_es_ready_0),
    .up_rdata_out (up_es_rdata_0_s),
    .up_ready_out (up_es_ready_0_s));

  assign up_ch_rst_0 = up_ch_rst;
  assign up_ch_user_ready_0 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_0 = up_ch_lpm_dfe_n;
  assign up_ch_rate_0 = up_ch_rate;
  assign up_ch_sys_clk_sel_0 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_0 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (0),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_0 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (1'd1),
    .up_rst_done_in (1'd1),
    .up_pll_locked (up_ch_pll_locked_0),
    .up_rst_done (up_ch_rst_done_0),
    .up_pll_locked_out (up_ch_pll_locked_0_s),
    .up_rst_done_out (up_ch_rst_done_0_s));

  assign up_ch_sel_0 = up_ch_sel;
  assign up_ch_enb_0 = up_ch_enb;
  assign up_ch_addr_0 = up_ch_addr;
  assign up_ch_wr_0 = up_ch_wr;
  assign up_ch_wdata_0 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (0),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_0 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (16'd0),
    .up_ready_in (1'd1),
    .up_rdata (up_ch_rdata_0),
    .up_ready (up_ch_ready_0),
    .up_rdata_out (up_ch_rdata_0_s),
    .up_ready_out (up_ch_ready_0_s));

  assign up_es_sel_1 = up_es_sel;
  assign up_es_enb_1 = up_es_enb;
  assign up_es_addr_1 = up_es_addr;
  assign up_es_wr_1 = up_es_wr;
  assign up_es_wdata_1 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (1),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_1 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_0_s),
    .up_ready_in (up_es_ready_0_s),
    .up_rdata (up_es_rdata_1),
    .up_ready (up_es_ready_1),
    .up_rdata_out (up_es_rdata_1_s),
    .up_ready_out (up_es_ready_1_s));

  assign up_ch_rst_1 = up_ch_rst;
  assign up_ch_user_ready_1 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_1 = up_ch_lpm_dfe_n;
  assign up_ch_rate_1 = up_ch_rate;
  assign up_ch_sys_clk_sel_1 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_1 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (1),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_1 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_0_s),
    .up_rst_done_in (up_ch_rst_done_0_s),
    .up_pll_locked (up_ch_pll_locked_1),
    .up_rst_done (up_ch_rst_done_1),
    .up_pll_locked_out (up_ch_pll_locked_1_s),
    .up_rst_done_out (up_ch_rst_done_1_s));

  assign up_ch_sel_1 = up_ch_sel;
  assign up_ch_enb_1 = up_ch_enb;
  assign up_ch_addr_1 = up_ch_addr;
  assign up_ch_wr_1 = up_ch_wr;
  assign up_ch_wdata_1 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (1),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_1 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_0_s),
    .up_ready_in (up_ch_ready_0_s),
    .up_rdata (up_ch_rdata_1),
    .up_ready (up_ch_ready_1),
    .up_rdata_out (up_ch_rdata_1_s),
    .up_ready_out (up_ch_ready_1_s));

  assign up_es_sel_2 = up_es_sel;
  assign up_es_enb_2 = up_es_enb;
  assign up_es_addr_2 = up_es_addr;
  assign up_es_wr_2 = up_es_wr;
  assign up_es_wdata_2 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (2),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_2 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_1_s),
    .up_ready_in (up_es_ready_1_s),
    .up_rdata (up_es_rdata_2),
    .up_ready (up_es_ready_2),
    .up_rdata_out (up_es_rdata_2_s),
    .up_ready_out (up_es_ready_2_s));

  assign up_ch_rst_2 = up_ch_rst;
  assign up_ch_user_ready_2 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_2 = up_ch_lpm_dfe_n;
  assign up_ch_rate_2 = up_ch_rate;
  assign up_ch_sys_clk_sel_2 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_2 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (2),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_2 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_1_s),
    .up_rst_done_in (up_ch_rst_done_1_s),
    .up_pll_locked (up_ch_pll_locked_2),
    .up_rst_done (up_ch_rst_done_2),
    .up_pll_locked_out (up_ch_pll_locked_2_s),
    .up_rst_done_out (up_ch_rst_done_2_s));

  assign up_ch_sel_2 = up_ch_sel;
  assign up_ch_enb_2 = up_ch_enb;
  assign up_ch_addr_2 = up_ch_addr;
  assign up_ch_wr_2 = up_ch_wr;
  assign up_ch_wdata_2 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (2),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_2 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_1_s),
    .up_ready_in (up_ch_ready_1_s),
    .up_rdata (up_ch_rdata_2),
    .up_ready (up_ch_ready_2),
    .up_rdata_out (up_ch_rdata_2_s),
    .up_ready_out (up_ch_ready_2_s));

  assign up_es_sel_3 = up_es_sel;
  assign up_es_enb_3 = up_es_enb;
  assign up_es_addr_3 = up_es_addr;
  assign up_es_wr_3 = up_es_wr;
  assign up_es_wdata_3 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (3),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_3 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_2_s),
    .up_ready_in (up_es_ready_2_s),
    .up_rdata (up_es_rdata_3),
    .up_ready (up_es_ready_3),
    .up_rdata_out (up_es_rdata_3_s),
    .up_ready_out (up_es_ready_3_s));

  assign up_ch_rst_3 = up_ch_rst;
  assign up_ch_user_ready_3 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_3 = up_ch_lpm_dfe_n;
  assign up_ch_rate_3 = up_ch_rate;
  assign up_ch_sys_clk_sel_3 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_3 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (3),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_3 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_2_s),
    .up_rst_done_in (up_ch_rst_done_2_s),
    .up_pll_locked (up_ch_pll_locked_3),
    .up_rst_done (up_ch_rst_done_3),
    .up_pll_locked_out (up_ch_pll_locked_3_s),
    .up_rst_done_out (up_ch_rst_done_3_s));

  assign up_ch_sel_3 = up_ch_sel;
  assign up_ch_enb_3 = up_ch_enb;
  assign up_ch_addr_3 = up_ch_addr;
  assign up_ch_wr_3 = up_ch_wr;
  assign up_ch_wdata_3 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (3),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_3 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_2_s),
    .up_ready_in (up_ch_ready_2_s),
    .up_rdata (up_ch_rdata_3),
    .up_ready (up_ch_ready_3),
    .up_rdata_out (up_ch_rdata_3_s),
    .up_ready_out (up_ch_ready_3_s));

  assign up_cm_sel_4 = up_cm_sel;
  assign up_cm_enb_4 = up_cm_enb;
  assign up_cm_addr_4 = up_cm_addr;
  assign up_cm_wr_4 = up_cm_wr;
  assign up_cm_wdata_4 = up_cm_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (4),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_cm_4 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_cm_sel),
    .up_enb (up_cm_enb),
    .up_rdata_in (up_cm_rdata_0_s),
    .up_ready_in (up_cm_ready_0_s),
    .up_rdata (up_cm_rdata_4),
    .up_ready (up_cm_ready_4),
    .up_rdata_out (up_cm_rdata_4_s),
    .up_ready_out (up_cm_ready_4_s));

  assign up_es_sel_4 = up_es_sel;
  assign up_es_enb_4 = up_es_enb;
  assign up_es_addr_4 = up_es_addr;
  assign up_es_wr_4 = up_es_wr;
  assign up_es_wdata_4 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (4),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_4 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_3_s),
    .up_ready_in (up_es_ready_3_s),
    .up_rdata (up_es_rdata_4),
    .up_ready (up_es_ready_4),
    .up_rdata_out (up_es_rdata_4_s),
    .up_ready_out (up_es_ready_4_s));

  assign up_ch_rst_4 = up_ch_rst;
  assign up_ch_user_ready_4 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_4 = up_ch_lpm_dfe_n;
  assign up_ch_rate_4 = up_ch_rate;
  assign up_ch_sys_clk_sel_4 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_4 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (4),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_4 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_3_s),
    .up_rst_done_in (up_ch_rst_done_3_s),
    .up_pll_locked (up_ch_pll_locked_4),
    .up_rst_done (up_ch_rst_done_4),
    .up_pll_locked_out (up_ch_pll_locked_4_s),
    .up_rst_done_out (up_ch_rst_done_4_s));

  assign up_ch_sel_4 = up_ch_sel;
  assign up_ch_enb_4 = up_ch_enb;
  assign up_ch_addr_4 = up_ch_addr;
  assign up_ch_wr_4 = up_ch_wr;
  assign up_ch_wdata_4 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (4),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_4 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_3_s),
    .up_ready_in (up_ch_ready_3_s),
    .up_rdata (up_ch_rdata_4),
    .up_ready (up_ch_ready_4),
    .up_rdata_out (up_ch_rdata_4_s),
    .up_ready_out (up_ch_ready_4_s));

  assign up_es_sel_5 = up_es_sel;
  assign up_es_enb_5 = up_es_enb;
  assign up_es_addr_5 = up_es_addr;
  assign up_es_wr_5 = up_es_wr;
  assign up_es_wdata_5 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (5),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_5 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_4_s),
    .up_ready_in (up_es_ready_4_s),
    .up_rdata (up_es_rdata_5),
    .up_ready (up_es_ready_5),
    .up_rdata_out (up_es_rdata_5_s),
    .up_ready_out (up_es_ready_5_s));

  assign up_ch_rst_5 = up_ch_rst;
  assign up_ch_user_ready_5 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_5 = up_ch_lpm_dfe_n;
  assign up_ch_rate_5 = up_ch_rate;
  assign up_ch_sys_clk_sel_5 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_5 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (5),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_5 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_4_s),
    .up_rst_done_in (up_ch_rst_done_4_s),
    .up_pll_locked (up_ch_pll_locked_5),
    .up_rst_done (up_ch_rst_done_5),
    .up_pll_locked_out (up_ch_pll_locked_5_s),
    .up_rst_done_out (up_ch_rst_done_5_s));

  assign up_ch_sel_5 = up_ch_sel;
  assign up_ch_enb_5 = up_ch_enb;
  assign up_ch_addr_5 = up_ch_addr;
  assign up_ch_wr_5 = up_ch_wr;
  assign up_ch_wdata_5 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (5),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_5 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_4_s),
    .up_ready_in (up_ch_ready_4_s),
    .up_rdata (up_ch_rdata_5),
    .up_ready (up_ch_ready_5),
    .up_rdata_out (up_ch_rdata_5_s),
    .up_ready_out (up_ch_ready_5_s));

  assign up_es_sel_6 = up_es_sel;
  assign up_es_enb_6 = up_es_enb;
  assign up_es_addr_6 = up_es_addr;
  assign up_es_wr_6 = up_es_wr;
  assign up_es_wdata_6 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (6),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_6 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_5_s),
    .up_ready_in (up_es_ready_5_s),
    .up_rdata (up_es_rdata_6),
    .up_ready (up_es_ready_6),
    .up_rdata_out (up_es_rdata_6_s),
    .up_ready_out (up_es_ready_6_s));

  assign up_ch_rst_6 = up_ch_rst;
  assign up_ch_user_ready_6 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_6 = up_ch_lpm_dfe_n;
  assign up_ch_rate_6 = up_ch_rate;
  assign up_ch_sys_clk_sel_6 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_6 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (6),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_6 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_5_s),
    .up_rst_done_in (up_ch_rst_done_5_s),
    .up_pll_locked (up_ch_pll_locked_6),
    .up_rst_done (up_ch_rst_done_6),
    .up_pll_locked_out (up_ch_pll_locked_6_s),
    .up_rst_done_out (up_ch_rst_done_6_s));

  assign up_ch_sel_6 = up_ch_sel;
  assign up_ch_enb_6 = up_ch_enb;
  assign up_ch_addr_6 = up_ch_addr;
  assign up_ch_wr_6 = up_ch_wr;
  assign up_ch_wdata_6 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (6),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_6 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_5_s),
    .up_ready_in (up_ch_ready_5_s),
    .up_rdata (up_ch_rdata_6),
    .up_ready (up_ch_ready_6),
    .up_rdata_out (up_ch_rdata_6_s),
    .up_ready_out (up_ch_ready_6_s));

  assign up_es_sel_7 = up_es_sel;
  assign up_es_enb_7 = up_es_enb;
  assign up_es_addr_7 = up_es_addr;
  assign up_es_wr_7 = up_es_wr;
  assign up_es_wdata_7 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (7),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_7 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_6_s),
    .up_ready_in (up_es_ready_6_s),
    .up_rdata (up_es_rdata_7),
    .up_ready (up_es_ready_7),
    .up_rdata_out (up_es_rdata_7_s),
    .up_ready_out (up_es_ready_7_s));

  assign up_ch_rst_7 = up_ch_rst;
  assign up_ch_user_ready_7 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_7 = up_ch_lpm_dfe_n;
  assign up_ch_rate_7 = up_ch_rate;
  assign up_ch_sys_clk_sel_7 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_7 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (7),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_7 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_6_s),
    .up_rst_done_in (up_ch_rst_done_6_s),
    .up_pll_locked (up_ch_pll_locked_7),
    .up_rst_done (up_ch_rst_done_7),
    .up_pll_locked_out (up_ch_pll_locked_7_s),
    .up_rst_done_out (up_ch_rst_done_7_s));

  assign up_ch_sel_7 = up_ch_sel;
  assign up_ch_enb_7 = up_ch_enb;
  assign up_ch_addr_7 = up_ch_addr;
  assign up_ch_wr_7 = up_ch_wr;
  assign up_ch_wdata_7 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (7),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_7 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_6_s),
    .up_ready_in (up_ch_ready_6_s),
    .up_rdata (up_ch_rdata_7),
    .up_ready (up_ch_ready_7),
    .up_rdata_out (up_ch_rdata_7_s),
    .up_ready_out (up_ch_ready_7_s));

  assign up_cm_sel_8 = up_cm_sel;
  assign up_cm_enb_8 = up_cm_enb;
  assign up_cm_addr_8 = up_cm_addr;
  assign up_cm_wr_8 = up_cm_wr;
  assign up_cm_wdata_8 = up_cm_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (8),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_cm_8 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_cm_sel),
    .up_enb (up_cm_enb),
    .up_rdata_in (up_cm_rdata_4_s),
    .up_ready_in (up_cm_ready_4_s),
    .up_rdata (up_cm_rdata_8),
    .up_ready (up_cm_ready_8),
    .up_rdata_out (up_cm_rdata_8_s),
    .up_ready_out (up_cm_ready_8_s));

  assign up_es_sel_8 = up_es_sel;
  assign up_es_enb_8 = up_es_enb;
  assign up_es_addr_8 = up_es_addr;
  assign up_es_wr_8 = up_es_wr;
  assign up_es_wdata_8 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (8),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_8 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_7_s),
    .up_ready_in (up_es_ready_7_s),
    .up_rdata (up_es_rdata_8),
    .up_ready (up_es_ready_8),
    .up_rdata_out (up_es_rdata_8_s),
    .up_ready_out (up_es_ready_8_s));

  assign up_ch_rst_8 = up_ch_rst;
  assign up_ch_user_ready_8 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_8 = up_ch_lpm_dfe_n;
  assign up_ch_rate_8 = up_ch_rate;
  assign up_ch_sys_clk_sel_8 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_8 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (8),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_8 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_7_s),
    .up_rst_done_in (up_ch_rst_done_7_s),
    .up_pll_locked (up_ch_pll_locked_8),
    .up_rst_done (up_ch_rst_done_8),
    .up_pll_locked_out (up_ch_pll_locked_8_s),
    .up_rst_done_out (up_ch_rst_done_8_s));

  assign up_ch_sel_8 = up_ch_sel;
  assign up_ch_enb_8 = up_ch_enb;
  assign up_ch_addr_8 = up_ch_addr;
  assign up_ch_wr_8 = up_ch_wr;
  assign up_ch_wdata_8 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (8),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_8 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_7_s),
    .up_ready_in (up_ch_ready_7_s),
    .up_rdata (up_ch_rdata_8),
    .up_ready (up_ch_ready_8),
    .up_rdata_out (up_ch_rdata_8_s),
    .up_ready_out (up_ch_ready_8_s));

  assign up_es_sel_9 = up_es_sel;
  assign up_es_enb_9 = up_es_enb;
  assign up_es_addr_9 = up_es_addr;
  assign up_es_wr_9 = up_es_wr;
  assign up_es_wdata_9 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (9),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_9 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_8_s),
    .up_ready_in (up_es_ready_8_s),
    .up_rdata (up_es_rdata_9),
    .up_ready (up_es_ready_9),
    .up_rdata_out (up_es_rdata_9_s),
    .up_ready_out (up_es_ready_9_s));

  assign up_ch_rst_9 = up_ch_rst;
  assign up_ch_user_ready_9 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_9 = up_ch_lpm_dfe_n;
  assign up_ch_rate_9 = up_ch_rate;
  assign up_ch_sys_clk_sel_9 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_9 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (9),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_9 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_8_s),
    .up_rst_done_in (up_ch_rst_done_8_s),
    .up_pll_locked (up_ch_pll_locked_9),
    .up_rst_done (up_ch_rst_done_9),
    .up_pll_locked_out (up_ch_pll_locked_9_s),
    .up_rst_done_out (up_ch_rst_done_9_s));

  assign up_ch_sel_9 = up_ch_sel;
  assign up_ch_enb_9 = up_ch_enb;
  assign up_ch_addr_9 = up_ch_addr;
  assign up_ch_wr_9 = up_ch_wr;
  assign up_ch_wdata_9 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (9),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_9 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_8_s),
    .up_ready_in (up_ch_ready_8_s),
    .up_rdata (up_ch_rdata_9),
    .up_ready (up_ch_ready_9),
    .up_rdata_out (up_ch_rdata_9_s),
    .up_ready_out (up_ch_ready_9_s));

  assign up_es_sel_10 = up_es_sel;
  assign up_es_enb_10 = up_es_enb;
  assign up_es_addr_10 = up_es_addr;
  assign up_es_wr_10 = up_es_wr;
  assign up_es_wdata_10 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (10),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_10 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_9_s),
    .up_ready_in (up_es_ready_9_s),
    .up_rdata (up_es_rdata_10),
    .up_ready (up_es_ready_10),
    .up_rdata_out (up_es_rdata_10_s),
    .up_ready_out (up_es_ready_10_s));

  assign up_ch_rst_10 = up_ch_rst;
  assign up_ch_user_ready_10 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_10 = up_ch_lpm_dfe_n;
  assign up_ch_rate_10 = up_ch_rate;
  assign up_ch_sys_clk_sel_10 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_10 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (10),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_10 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_9_s),
    .up_rst_done_in (up_ch_rst_done_9_s),
    .up_pll_locked (up_ch_pll_locked_10),
    .up_rst_done (up_ch_rst_done_10),
    .up_pll_locked_out (up_ch_pll_locked_10_s),
    .up_rst_done_out (up_ch_rst_done_10_s));

  assign up_ch_sel_10 = up_ch_sel;
  assign up_ch_enb_10 = up_ch_enb;
  assign up_ch_addr_10 = up_ch_addr;
  assign up_ch_wr_10 = up_ch_wr;
  assign up_ch_wdata_10 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (10),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_10 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_9_s),
    .up_ready_in (up_ch_ready_9_s),
    .up_rdata (up_ch_rdata_10),
    .up_ready (up_ch_ready_10),
    .up_rdata_out (up_ch_rdata_10_s),
    .up_ready_out (up_ch_ready_10_s));

  assign up_es_sel_11 = up_es_sel;
  assign up_es_enb_11 = up_es_enb;
  assign up_es_addr_11 = up_es_addr;
  assign up_es_wr_11 = up_es_wr;
  assign up_es_wdata_11 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (11),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_11 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_10_s),
    .up_ready_in (up_es_ready_10_s),
    .up_rdata (up_es_rdata_11),
    .up_ready (up_es_ready_11),
    .up_rdata_out (up_es_rdata_11_s),
    .up_ready_out (up_es_ready_11_s));

  assign up_ch_rst_11 = up_ch_rst;
  assign up_ch_user_ready_11 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_11 = up_ch_lpm_dfe_n;
  assign up_ch_rate_11 = up_ch_rate;
  assign up_ch_sys_clk_sel_11 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_11 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (11),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_11 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_10_s),
    .up_rst_done_in (up_ch_rst_done_10_s),
    .up_pll_locked (up_ch_pll_locked_11),
    .up_rst_done (up_ch_rst_done_11),
    .up_pll_locked_out (up_ch_pll_locked_11_s),
    .up_rst_done_out (up_ch_rst_done_11_s));

  assign up_ch_sel_11 = up_ch_sel;
  assign up_ch_enb_11 = up_ch_enb;
  assign up_ch_addr_11 = up_ch_addr;
  assign up_ch_wr_11 = up_ch_wr;
  assign up_ch_wdata_11 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (11),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_11 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_10_s),
    .up_ready_in (up_ch_ready_10_s),
    .up_rdata (up_ch_rdata_11),
    .up_ready (up_ch_ready_11),
    .up_rdata_out (up_ch_rdata_11_s),
    .up_ready_out (up_ch_ready_11_s));

  assign up_cm_sel_12 = up_cm_sel;
  assign up_cm_enb_12 = up_cm_enb;
  assign up_cm_addr_12 = up_cm_addr;
  assign up_cm_wr_12 = up_cm_wr;
  assign up_cm_wdata_12 = up_cm_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (12),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_cm_12 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_cm_sel),
    .up_enb (up_cm_enb),
    .up_rdata_in (up_cm_rdata_8_s),
    .up_ready_in (up_cm_ready_8_s),
    .up_rdata (up_cm_rdata_12),
    .up_ready (up_cm_ready_12),
    .up_rdata_out (up_cm_rdata_12_s),
    .up_ready_out (up_cm_ready_12_s));

  assign up_es_sel_12 = up_es_sel;
  assign up_es_enb_12 = up_es_enb;
  assign up_es_addr_12 = up_es_addr;
  assign up_es_wr_12 = up_es_wr;
  assign up_es_wdata_12 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (12),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_12 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_11_s),
    .up_ready_in (up_es_ready_11_s),
    .up_rdata (up_es_rdata_12),
    .up_ready (up_es_ready_12),
    .up_rdata_out (up_es_rdata_12_s),
    .up_ready_out (up_es_ready_12_s));

  assign up_ch_rst_12 = up_ch_rst;
  assign up_ch_user_ready_12 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_12 = up_ch_lpm_dfe_n;
  assign up_ch_rate_12 = up_ch_rate;
  assign up_ch_sys_clk_sel_12 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_12 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (12),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_12 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_11_s),
    .up_rst_done_in (up_ch_rst_done_11_s),
    .up_pll_locked (up_ch_pll_locked_12),
    .up_rst_done (up_ch_rst_done_12),
    .up_pll_locked_out (up_ch_pll_locked_12_s),
    .up_rst_done_out (up_ch_rst_done_12_s));

  assign up_ch_sel_12 = up_ch_sel;
  assign up_ch_enb_12 = up_ch_enb;
  assign up_ch_addr_12 = up_ch_addr;
  assign up_ch_wr_12 = up_ch_wr;
  assign up_ch_wdata_12 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (12),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_12 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_11_s),
    .up_ready_in (up_ch_ready_11_s),
    .up_rdata (up_ch_rdata_12),
    .up_ready (up_ch_ready_12),
    .up_rdata_out (up_ch_rdata_12_s),
    .up_ready_out (up_ch_ready_12_s));

  assign up_es_sel_13 = up_es_sel;
  assign up_es_enb_13 = up_es_enb;
  assign up_es_addr_13 = up_es_addr;
  assign up_es_wr_13 = up_es_wr;
  assign up_es_wdata_13 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (13),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_13 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_12_s),
    .up_ready_in (up_es_ready_12_s),
    .up_rdata (up_es_rdata_13),
    .up_ready (up_es_ready_13),
    .up_rdata_out (up_es_rdata_13_s),
    .up_ready_out (up_es_ready_13_s));

  assign up_ch_rst_13 = up_ch_rst;
  assign up_ch_user_ready_13 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_13 = up_ch_lpm_dfe_n;
  assign up_ch_rate_13 = up_ch_rate;
  assign up_ch_sys_clk_sel_13 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_13 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (13),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_13 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_12_s),
    .up_rst_done_in (up_ch_rst_done_12_s),
    .up_pll_locked (up_ch_pll_locked_13),
    .up_rst_done (up_ch_rst_done_13),
    .up_pll_locked_out (up_ch_pll_locked_13_s),
    .up_rst_done_out (up_ch_rst_done_13_s));

  assign up_ch_sel_13 = up_ch_sel;
  assign up_ch_enb_13 = up_ch_enb;
  assign up_ch_addr_13 = up_ch_addr;
  assign up_ch_wr_13 = up_ch_wr;
  assign up_ch_wdata_13 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (13),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_13 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_12_s),
    .up_ready_in (up_ch_ready_12_s),
    .up_rdata (up_ch_rdata_13),
    .up_ready (up_ch_ready_13),
    .up_rdata_out (up_ch_rdata_13_s),
    .up_ready_out (up_ch_ready_13_s));

  assign up_es_sel_14 = up_es_sel;
  assign up_es_enb_14 = up_es_enb;
  assign up_es_addr_14 = up_es_addr;
  assign up_es_wr_14 = up_es_wr;
  assign up_es_wdata_14 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (14),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_14 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_13_s),
    .up_ready_in (up_es_ready_13_s),
    .up_rdata (up_es_rdata_14),
    .up_ready (up_es_ready_14),
    .up_rdata_out (up_es_rdata_14_s),
    .up_ready_out (up_es_ready_14_s));

  assign up_ch_rst_14 = up_ch_rst;
  assign up_ch_user_ready_14 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_14 = up_ch_lpm_dfe_n;
  assign up_ch_rate_14 = up_ch_rate;
  assign up_ch_sys_clk_sel_14 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_14 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (14),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_14 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_13_s),
    .up_rst_done_in (up_ch_rst_done_13_s),
    .up_pll_locked (up_ch_pll_locked_14),
    .up_rst_done (up_ch_rst_done_14),
    .up_pll_locked_out (up_ch_pll_locked_14_s),
    .up_rst_done_out (up_ch_rst_done_14_s));

  assign up_ch_sel_14 = up_ch_sel;
  assign up_ch_enb_14 = up_ch_enb;
  assign up_ch_addr_14 = up_ch_addr;
  assign up_ch_wr_14 = up_ch_wr;
  assign up_ch_wdata_14 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (14),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_14 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_13_s),
    .up_ready_in (up_ch_ready_13_s),
    .up_rdata (up_ch_rdata_14),
    .up_ready (up_ch_ready_14),
    .up_rdata_out (up_ch_rdata_14_s),
    .up_ready_out (up_ch_ready_14_s));

  assign up_es_sel_15 = up_es_sel;
  assign up_es_enb_15 = up_es_enb;
  assign up_es_addr_15 = up_es_addr;
  assign up_es_wr_15 = up_es_wr;
  assign up_es_wdata_15 = up_es_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (15),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_es_15 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_es_sel),
    .up_enb (up_es_enb),
    .up_rdata_in (up_es_rdata_14_s),
    .up_ready_in (up_es_ready_14_s),
    .up_rdata (up_es_rdata_15),
    .up_ready (up_es_ready_15),
    .up_rdata_out (up_es_rdata_15_s),
    .up_ready_out (up_es_ready_15_s));

  assign up_ch_rst_15 = up_ch_rst;
  assign up_ch_user_ready_15 = up_ch_user_ready;
  assign up_ch_lpm_dfe_n_15 = up_ch_lpm_dfe_n;
  assign up_ch_rate_15 = up_ch_rate;
  assign up_ch_sys_clk_sel_15 = up_ch_sys_clk_sel;
  assign up_ch_out_clk_sel_15 = up_ch_out_clk_sel;

  axi_adxcvr_mstatus #(
    .XCVR_ID (15),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mstatus_ch_15 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_pll_locked_in (up_ch_pll_locked_14_s),
    .up_rst_done_in (up_ch_rst_done_14_s),
    .up_pll_locked (up_ch_pll_locked_15),
    .up_rst_done (up_ch_rst_done_15),
    .up_pll_locked_out (up_ch_pll_locked_15_s),
    .up_rst_done_out (up_ch_rst_done_15_s));

  assign up_ch_sel_15 = up_ch_sel;
  assign up_ch_enb_15 = up_ch_enb;
  assign up_ch_addr_15 = up_ch_addr;
  assign up_ch_wr_15 = up_ch_wr;
  assign up_ch_wdata_15 = up_ch_wdata;

  axi_adxcvr_mdrp #(
    .XCVR_ID (15),
    .NUM_OF_LANES (NUM_OF_LANES))
  i_mdrp_ch_15 (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_sel (up_ch_sel),
    .up_enb (up_ch_enb),
    .up_rdata_in (up_ch_rdata_14_s),
    .up_ready_in (up_ch_ready_14_s),
    .up_rdata (up_ch_rdata_15),
    .up_ready (up_ch_ready_15),
    .up_rdata_out (up_ch_rdata_15_s),
    .up_ready_out (up_ch_ready_15_s));

  axi_adxcvr_es #(
    .GTH_OR_GTX_N (GTH_OR_GTX_N),
    .TX_OR_RX_N (TX_OR_RX_N))
  i_es (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_es_enb (up_es_enb),
    .up_es_addr (up_es_addr),
    .up_es_wr (up_es_wr),
    .up_es_wdata (up_es_wdata),
    .up_es_rdata (up_es_rdata_15_s),
    .up_es_ready (up_es_ready_15_s),
    .up_ch_lpm_dfe_n (up_ch_lpm_dfe_n),
    .up_es_req (up_es_req),
    .up_es_ack (up_es_ack),
    .up_es_pscale (up_es_pscale),
    .up_es_vrange (up_es_vrange),
    .up_es_vstep (up_es_vstep),
    .up_es_vmax (up_es_vmax),
    .up_es_vmin (up_es_vmin),
    .up_es_hmax (up_es_hmax),
    .up_es_hmin (up_es_hmin),
    .up_es_hstep (up_es_hstep),
    .up_es_saddr (up_es_saddr),
    .up_es_status (up_es_status),
    .up_axi_awvalid (m_axi_awvalid),
    .up_axi_awaddr (m_axi_awaddr),
    .up_axi_awprot (m_axi_awprot),
    .up_axi_awready (m_axi_awready),
    .up_axi_wvalid (m_axi_wvalid),
    .up_axi_wdata (m_axi_wdata),
    .up_axi_wstrb (m_axi_wstrb),
    .up_axi_wready (m_axi_wready),
    .up_axi_bvalid (m_axi_bvalid),
    .up_axi_bresp (m_axi_bresp),
    .up_axi_bready (m_axi_bready),
    .up_axi_arvalid (m_axi_arvalid),
    .up_axi_araddr (m_axi_araddr),
    .up_axi_arprot (m_axi_arprot),
    .up_axi_arready (m_axi_arready),
    .up_axi_rvalid (m_axi_rvalid),
    .up_axi_rdata (m_axi_rdata),
    .up_axi_rresp (m_axi_rresp),
    .up_axi_rready (m_axi_rready));

  axi_adxcvr_up #(
    .ID (ID),
    .NUM_OF_LANES (NUM_OF_LANES),
    .GTH_OR_GTX_N (GTH_OR_GTX_N),
    .TX_OR_RX_N (TX_OR_RX_N),
    .QPLL_ENABLE (QPLL_ENABLE),
    .LPM_OR_DFE_N (LPM_OR_DFE_N),
    .RATE (RATE),
    .SYS_CLK_SEL (SYS_CLK_SEL),
    .OUT_CLK_SEL (OUT_CLK_SEL))
  i_up (
    .up_cm_sel (up_cm_sel),
    .up_cm_enb (up_cm_enb),
    .up_cm_addr (up_cm_addr),
    .up_cm_wr (up_cm_wr),
    .up_cm_wdata (up_cm_wdata),
    .up_cm_rdata (up_cm_rdata_12_s),
    .up_cm_ready (up_cm_ready_12_s),
    .up_ch_pll_locked (up_ch_pll_locked_15_s),
    .up_ch_rst (up_ch_rst),
    .up_ch_user_ready (up_ch_user_ready),
    .up_ch_rst_done (up_ch_rst_done_15_s),
    .up_ch_lpm_dfe_n (up_ch_lpm_dfe_n),
    .up_ch_rate (up_ch_rate),
    .up_ch_sys_clk_sel (up_ch_sys_clk_sel),
    .up_ch_out_clk_sel (up_ch_out_clk_sel),
    .up_ch_sel (up_ch_sel),
    .up_ch_enb (up_ch_enb),
    .up_ch_addr (up_ch_addr),
    .up_ch_wr (up_ch_wr),
    .up_ch_wdata (up_ch_wdata),
    .up_ch_rdata (up_ch_rdata_15_s),
    .up_ch_ready (up_ch_ready_15_s),
    .up_es_sel (up_es_sel),
    .up_es_req (up_es_req),
    .up_es_ack (up_es_ack),
    .up_es_pscale (up_es_pscale),
    .up_es_vrange (up_es_vrange),
    .up_es_vstep (up_es_vstep),
    .up_es_vmax (up_es_vmax),
    .up_es_vmin (up_es_vmin),
    .up_es_hmax (up_es_hmax),
    .up_es_hmin (up_es_hmin),
    .up_es_hstep (up_es_hstep),
    .up_es_saddr (up_es_saddr),
    .up_es_status (up_es_status),
    .up_status (up_status),
    .up_pll_rst (up_pll_rst),
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_wreq (up_wreq),
    .up_waddr (up_waddr),
    .up_wdata (up_wdata),
    .up_wack (up_wack),
    .up_rreq (up_rreq),
    .up_raddr (up_raddr),
    .up_rdata (up_rdata),
    .up_rack (up_rack));

  up_axi #(.ADDRESS_WIDTH (10)) i_axi (
    .up_rstn (up_rstn),
    .up_clk (up_clk),
    .up_axi_awvalid (s_axi_awvalid),
    .up_axi_awaddr (s_axi_awaddr),
    .up_axi_awready (s_axi_awready),
    .up_axi_wvalid (s_axi_wvalid),
    .up_axi_wdata (s_axi_wdata),
    .up_axi_wstrb (s_axi_wstrb),
    .up_axi_wready (s_axi_wready),
    .up_axi_bvalid (s_axi_bvalid),
    .up_axi_bresp (s_axi_bresp),
    .up_axi_bready (s_axi_bready),
    .up_axi_arvalid (s_axi_arvalid),
    .up_axi_araddr (s_axi_araddr),
    .up_axi_arready (s_axi_arready),
    .up_axi_rvalid (s_axi_rvalid),
    .up_axi_rresp (s_axi_rresp),
    .up_axi_rdata (s_axi_rdata),
    .up_axi_rready (s_axi_rready),
    .up_wreq (up_wreq),
    .up_waddr (up_waddr),
    .up_wdata (up_wdata),
    .up_wack (up_wack),
    .up_rreq (up_rreq),
    .up_raddr (up_raddr),
    .up_rdata (up_rdata),
    .up_rack (up_rack));

endmodule

// ***************************************************************************
// ***************************************************************************

